/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu May  6 01:56:08 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 721959473 */

module datapath(B, A, Z);
   input [15:0]B;
   input [15:0]A;
   output [31:0]Z;

   HA_X1 i_0 (.A(n_262), .B(n_277), .CO(n_285), .S(n_284));
   FA_X1 i_1 (.A(n_272), .B(n_278), .CI(n_295), .CO(n_301), .S(n_300));
   HA_X1 i_2 (.A(n_288), .B(n_285), .CO(n_303), .S(n_302));
   FA_X1 i_3 (.A(n_313), .B(n_306), .CI(n_320), .CO(n_327), .S(n_326));
   HA_X1 i_4 (.A(n_303), .B(n_301), .CO(n_329), .S(n_328));
   FA_X1 i_5 (.A(n_307), .B(n_321), .CI(n_345), .CO(n_353), .S(n_352));
   FA_X1 i_6 (.A(n_339), .B(n_332), .CI(n_329), .CO(n_355), .S(n_354));
   HA_X1 i_7 (.A(n_352), .B(n_327), .CO(n_357), .S(n_356));
   FA_X1 i_8 (.A(n_340), .B(n_333), .CI(n_346), .CO(n_380), .S(n_379));
   FA_X1 i_9 (.A(n_374), .B(n_367), .CI(n_360), .CO(n_382), .S(n_381));
   FA_X1 i_10 (.A(n_379), .B(n_353), .CI(n_357), .CO(n_384), .S(n_383));
   HA_X1 i_11 (.A(n_355), .B(n_381), .CO(n_386), .S(n_385));
   FA_X1 i_12 (.A(n_361), .B(n_403), .CI(n_396), .CO(n_417), .S(n_416));
   FA_X1 i_13 (.A(n_389), .B(n_380), .CI(n_410), .CO(n_419), .S(n_418));
   FA_X1 i_14 (.A(n_382), .B(n_416), .CI(n_418), .CO(n_421), .S(n_420));
   HA_X1 i_15 (.A(n_386), .B(n_384), .CO(n_423), .S(n_422));
   FA_X1 i_16 (.A(n_397), .B(n_390), .CI(n_411), .CO(n_454), .S(n_453));
   FA_X1 i_17 (.A(n_446), .B(n_440), .CI(n_433), .CO(n_456), .S(n_455));
   FA_X1 i_18 (.A(n_426), .B(n_453), .CI(n_417), .CO(n_458), .S(n_457));
   FA_X1 i_19 (.A(n_419), .B(n_455), .CI(n_457), .CO(n_460), .S(n_459));
   HA_X1 i_20 (.A(n_423), .B(n_421), .CO(n_462), .S(n_461));
   FA_X1 i_21 (.A(n_441), .B(n_434), .CI(n_427), .CO(n_492), .S(n_491));
   FA_X1 i_22 (.A(n_447), .B(n_486), .CI(n_479), .CO(n_494), .S(n_493));
   FA_X1 i_23 (.A(n_472), .B(n_465), .CI(n_454), .CO(n_496), .S(n_495));
   FA_X1 i_24 (.A(n_491), .B(n_456), .CI(n_458), .CO(n_498), .S(n_497));
   FA_X1 i_25 (.A(n_495), .B(n_493), .CI(n_497), .CO(n_500), .S(n_499));
   HA_X1 i_26 (.A(n_462), .B(n_460), .CO(n_502), .S(n_501));
   FA_X1 i_27 (.A(n_473), .B(n_466), .CI(n_492), .CO(n_540), .S(n_539));
   FA_X1 i_28 (.A(n_526), .B(n_519), .CI(n_512), .CO(n_542), .S(n_541));
   FA_X1 i_29 (.A(n_505), .B(n_539), .CI(n_533), .CO(n_544), .S(n_543));
   FA_X1 i_30 (.A(n_494), .B(n_496), .CI(n_541), .CO(n_546), .S(n_545));
   FA_X1 i_31 (.A(n_498), .B(n_543), .CI(n_545), .CO(n_548), .S(n_547));
   HA_X1 i_32 (.A(n_500), .B(n_502), .CO(n_550), .S(n_549));
   FA_X1 i_33 (.A(n_520), .B(n_513), .CI(n_506), .CO(n_588), .S(n_587));
   FA_X1 i_34 (.A(n_534), .B(n_580), .CI(n_574), .CO(n_590), .S(n_589));
   FA_X1 i_35 (.A(n_567), .B(n_560), .CI(n_553), .CO(n_592), .S(n_591));
   FA_X1 i_36 (.A(n_540), .B(n_587), .CI(n_542), .CO(n_594), .S(n_593));
   FA_X1 i_37 (.A(n_544), .B(n_591), .CI(n_589), .CO(n_596), .S(n_595));
   FA_X1 i_38 (.A(n_593), .B(n_546), .CI(n_548), .CO(n_598), .S(n_597));
   HA_X1 i_39 (.A(n_595), .B(n_550), .CO(n_600), .S(n_599));
   FA_X1 i_40 (.A(n_575), .B(n_568), .CI(n_561), .CO(n_637), .S(n_636));
   FA_X1 i_41 (.A(n_554), .B(n_588), .CI(n_581), .CO(n_639), .S(n_638));
   FA_X1 i_42 (.A(n_631), .B(n_624), .CI(n_617), .CO(n_641), .S(n_640));
   FA_X1 i_43 (.A(n_610), .B(n_603), .CI(n_636), .CO(n_643), .S(n_642));
   FA_X1 i_44 (.A(n_592), .B(n_590), .CI(n_638), .CO(n_645), .S(n_644));
   FA_X1 i_45 (.A(n_594), .B(n_642), .CI(n_640), .CO(n_647), .S(n_646));
   FA_X1 i_46 (.A(n_644), .B(n_596), .CI(n_646), .CO(n_649), .S(n_648));
   HA_X1 i_47 (.A(n_598), .B(n_600), .CO(n_651), .S(n_650));
   FA_X1 i_48 (.A(n_618), .B(n_611), .CI(n_604), .CO(n_696), .S(n_695));
   FA_X1 i_49 (.A(n_637), .B(n_682), .CI(n_675), .CO(n_698), .S(n_697));
   FA_X1 i_50 (.A(n_668), .B(n_661), .CI(n_654), .CO(n_700), .S(n_699));
   FA_X1 i_51 (.A(n_639), .B(n_695), .CI(n_689), .CO(n_702), .S(n_701));
   FA_X1 i_52 (.A(n_641), .B(n_643), .CI(n_699), .CO(n_704), .S(n_703));
   FA_X1 i_53 (.A(n_697), .B(n_645), .CI(n_701), .CO(n_706), .S(n_705));
   FA_X1 i_54 (.A(n_647), .B(n_703), .CI(n_705), .CO(n_708), .S(n_707));
   HA_X1 i_55 (.A(n_649), .B(n_651), .CO(n_710), .S(n_709));
   FA_X1 i_56 (.A(n_683), .B(n_676), .CI(n_669), .CO(n_747), .S(n_746));
   FA_X1 i_57 (.A(n_662), .B(n_655), .CI(n_696), .CO(n_749), .S(n_748));
   FA_X1 i_58 (.A(n_690), .B(n_741), .CI(n_734), .CO(n_751), .S(n_750));
   FA_X1 i_59 (.A(n_727), .B(n_720), .CI(n_713), .CO(n_753), .S(n_752));
   FA_X1 i_60 (.A(n_748), .B(n_746), .CI(n_700), .CO(n_755), .S(n_754));
   FA_X1 i_61 (.A(n_698), .B(n_702), .CI(n_752), .CO(n_757), .S(n_756));
   FA_X1 i_62 (.A(n_750), .B(n_754), .CI(n_704), .CO(n_759), .S(n_758));
   FA_X1 i_63 (.A(n_756), .B(n_706), .CI(n_758), .CO(n_761), .S(n_760));
   HA_X1 i_64 (.A(n_708), .B(n_710), .CO(n_763), .S(n_762));
   FA_X1 i_65 (.A(n_735), .B(n_728), .CI(n_721), .CO(n_801), .S(n_800));
   FA_X1 i_66 (.A(n_714), .B(n_747), .CI(n_793), .CO(n_803), .S(n_802));
   FA_X1 i_67 (.A(n_787), .B(n_780), .CI(n_773), .CO(n_805), .S(n_804));
   FA_X1 i_68 (.A(n_766), .B(n_749), .CI(n_800), .CO(n_807), .S(n_806));
   FA_X1 i_69 (.A(n_753), .B(n_751), .CI(n_802), .CO(n_809), .S(n_808));
   FA_X1 i_70 (.A(n_755), .B(n_804), .CI(n_806), .CO(n_811), .S(n_810));
   FA_X1 i_71 (.A(n_808), .B(n_757), .CI(n_759), .CO(n_813), .S(n_812));
   FA_X1 i_72 (.A(n_810), .B(n_812), .CI(n_761), .CO(n_815), .S(n_814));
   FA_X1 i_73 (.A(n_774), .B(n_767), .CI(n_801), .CO(n_853), .S(n_852));
   FA_X1 i_74 (.A(n_794), .B(n_839), .CI(n_832), .CO(n_855), .S(n_854));
   FA_X1 i_75 (.A(n_825), .B(n_818), .CI(n_852), .CO(n_857), .S(n_856));
   FA_X1 i_76 (.A(n_846), .B(n_805), .CI(n_803), .CO(n_859), .S(n_858));
   FA_X1 i_77 (.A(n_807), .B(n_856), .CI(n_854), .CO(n_861), .S(n_860));
   FA_X1 i_78 (.A(n_809), .B(n_858), .CI(n_811), .CO(n_863), .S(n_862));
   FA_X1 i_79 (.A(n_860), .B(n_813), .CI(n_862), .CO(n_865), .S(n_864));
   FA_X1 i_80 (.A(n_840), .B(n_833), .CI(n_826), .CO(n_895), .S(n_894));
   FA_X1 i_81 (.A(n_819), .B(n_847), .CI(n_889), .CO(n_897), .S(n_896));
   FA_X1 i_82 (.A(n_882), .B(n_875), .CI(n_868), .CO(n_899), .S(n_898));
   FA_X1 i_83 (.A(n_853), .B(n_894), .CI(n_855), .CO(n_901), .S(n_900));
   FA_X1 i_84 (.A(n_896), .B(n_859), .CI(n_857), .CO(n_903), .S(n_902));
   FA_X1 i_85 (.A(n_898), .B(n_900), .CI(n_861), .CO(n_905), .S(n_904));
   FA_X1 i_86 (.A(n_902), .B(n_863), .CI(n_904), .CO(n_907), .S(n_906));
   FA_X1 i_87 (.A(n_883), .B(n_876), .CI(n_869), .CO(n_938), .S(n_937));
   FA_X1 i_88 (.A(n_895), .B(n_930), .CI(n_924), .CO(n_940), .S(n_939));
   FA_X1 i_89 (.A(n_917), .B(n_910), .CI(n_937), .CO(n_942), .S(n_941));
   FA_X1 i_90 (.A(n_899), .B(n_897), .CI(n_901), .CO(n_944), .S(n_943));
   FA_X1 i_91 (.A(n_941), .B(n_939), .CI(n_903), .CO(n_946), .S(n_945));
   FA_X1 i_92 (.A(n_943), .B(n_905), .CI(n_945), .CO(n_948), .S(n_947));
   FA_X1 i_93 (.A(n_911), .B(n_938), .CI(n_931), .CO(n_1), .S(n_0));
   FA_X1 i_94 (.A(n_105), .B(n_958), .CI(n_951), .CO(n_3), .S(n_2));
   FA_X1 i_95 (.A(n_104), .B(n_940), .CI(n_0), .CO(n_5), .S(n_4));
   FA_X1 i_96 (.A(n_942), .B(n_2), .CI(n_944), .CO(n_7), .S(n_6));
   FA_X1 i_97 (.A(n_4), .B(n_946), .CI(n_6), .CO(n_9), .S(n_8));
   FA_X1 i_98 (.A(n_103), .B(n_959), .CI(n_952), .CO(n_11), .S(n_10));
   FA_X1 i_99 (.A(n_102), .B(n_101), .CI(n_100), .CO(n_13), .S(n_12));
   FA_X1 i_100 (.A(n_99), .B(n_1), .CI(n_10), .CO(n_15), .S(n_14));
   FA_X1 i_101 (.A(n_3), .B(n_12), .CI(n_14), .CO(n_17), .S(n_16));
   FA_X1 i_102 (.A(n_5), .B(n_7), .CI(n_16), .CO(n_19), .S(n_18));
   FA_X1 i_103 (.A(n_98), .B(n_97), .CI(n_11), .CO(n_21), .S(n_20));
   FA_X1 i_104 (.A(n_96), .B(n_95), .CI(n_94), .CO(n_23), .S(n_22));
   FA_X1 i_105 (.A(n_20), .B(n_13), .CI(n_15), .CO(n_25), .S(n_24));
   FA_X1 i_106 (.A(n_22), .B(n_24), .CI(n_17), .CO(n_27), .S(n_26));
   FA_X1 i_107 (.A(n_93), .B(n_92), .CI(n_91), .CO(n_29), .S(n_28));
   FA_X1 i_108 (.A(n_21), .B(n_90), .CI(n_23), .CO(n_31), .S(n_30));
   FA_X1 i_109 (.A(n_28), .B(n_25), .CI(n_30), .CO(n_33), .S(n_32));
   FA_X1 i_110 (.A(n_89), .B(n_88), .CI(n_87), .CO(n_35), .S(n_34));
   FA_X1 i_111 (.A(n_86), .B(n_85), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_112 (.A(n_29), .B(n_31), .CI(n_36), .CO(n_39), .S(n_38));
   FA_X1 i_113 (.A(n_84), .B(n_83), .CI(n_82), .CO(n_41), .S(n_40));
   FA_X1 i_114 (.A(n_35), .B(n_37), .CI(n_40), .CO(n_43), .S(n_42));
   FA_X1 i_115 (.A(n_81), .B(n_80), .CI(n_41), .CO(n_45), .S(n_44));
   FA_X1 i_116 (.A(n_79), .B(n_78), .CI(n_77), .CO(n_47), .S(n_46));
   FA_X1 i_117 (.A(n_266), .B(n_261), .CI(n_76), .CO(n_48), .S(Z[3]));
   FA_X1 i_118 (.A(n_271), .B(n_284), .CI(n_48), .CO(n_49), .S(Z[4]));
   FA_X1 i_119 (.A(n_302), .B(n_300), .CI(n_49), .CO(n_50), .S(Z[5]));
   FA_X1 i_120 (.A(n_328), .B(n_326), .CI(n_50), .CO(n_51), .S(Z[6]));
   FA_X1 i_121 (.A(n_354), .B(n_356), .CI(n_51), .CO(n_52), .S(Z[7]));
   FA_X1 i_122 (.A(n_383), .B(n_385), .CI(n_52), .CO(n_53), .S(Z[8]));
   FA_X1 i_123 (.A(n_422), .B(n_420), .CI(n_53), .CO(n_54), .S(Z[9]));
   FA_X1 i_124 (.A(n_461), .B(n_459), .CI(n_54), .CO(n_55), .S(Z[10]));
   FA_X1 i_125 (.A(n_499), .B(n_501), .CI(n_55), .CO(n_56), .S(Z[11]));
   FA_X1 i_126 (.A(n_547), .B(n_549), .CI(n_56), .CO(n_57), .S(Z[12]));
   FA_X1 i_127 (.A(n_597), .B(n_599), .CI(n_57), .CO(n_58), .S(Z[13]));
   FA_X1 i_128 (.A(n_648), .B(n_650), .CI(n_58), .CO(n_59), .S(Z[14]));
   FA_X1 i_129 (.A(n_707), .B(n_709), .CI(n_59), .CO(n_60), .S(Z[15]));
   FA_X1 i_130 (.A(n_760), .B(n_762), .CI(n_60), .CO(n_61), .S(Z[16]));
   FA_X1 i_131 (.A(n_763), .B(n_814), .CI(n_61), .CO(n_62), .S(Z[17]));
   FA_X1 i_132 (.A(n_864), .B(n_815), .CI(n_62), .CO(n_63), .S(Z[18]));
   FA_X1 i_133 (.A(n_865), .B(n_906), .CI(n_63), .CO(n_64), .S(Z[19]));
   FA_X1 i_134 (.A(n_947), .B(n_907), .CI(n_64), .CO(n_65), .S(Z[20]));
   FA_X1 i_135 (.A(n_948), .B(n_8), .CI(n_65), .CO(n_66), .S(Z[21]));
   FA_X1 i_136 (.A(n_9), .B(n_18), .CI(n_66), .CO(n_67), .S(Z[22]));
   FA_X1 i_137 (.A(n_26), .B(n_19), .CI(n_67), .CO(n_68), .S(Z[23]));
   FA_X1 i_138 (.A(n_27), .B(n_32), .CI(n_68), .CO(n_69), .S(Z[24]));
   FA_X1 i_139 (.A(n_38), .B(n_33), .CI(n_69), .CO(n_70), .S(Z[25]));
   FA_X1 i_140 (.A(n_39), .B(n_42), .CI(n_70), .CO(n_71), .S(Z[26]));
   FA_X1 i_141 (.A(n_44), .B(n_43), .CI(n_71), .CO(n_72), .S(Z[27]));
   FA_X1 i_142 (.A(n_45), .B(n_46), .CI(n_72), .CO(n_73), .S(Z[28]));
   FA_X1 i_143 (.A(n_75), .B(n_47), .CI(n_73), .CO(n_74), .S(Z[29]));
   NAND2_X1 i_144 (.A1(A[14]), .A2(B[14]), .ZN(n_106));
   INV_X1 i_145 (.A(n_106), .ZN(n_107));
   NAND3_X1 i_146 (.A1(n_107), .A2(B[15]), .A3(A[13]), .ZN(n_108));
   INV_X1 i_147 (.A(n_108), .ZN(n_109));
   INV_X1 i_148 (.A(B[15]), .ZN(n_110));
   INV_X1 i_149 (.A(A[13]), .ZN(n_111));
   OAI21_X1 i_150 (.A(n_106), .B1(n_110), .B2(n_111), .ZN(n_112));
   AND2_X1 i_151 (.A1(A[15]), .A2(B[13]), .ZN(n_113));
   AOI21_X1 i_152 (.A(n_109), .B1(n_112), .B2(n_113), .ZN(n_114));
   NAND2_X1 i_153 (.A1(A[15]), .A2(B[15]), .ZN(n_115));
   NOR2_X1 i_154 (.A1(n_106), .A2(n_115), .ZN(n_116));
   AOI22_X1 i_155 (.A1(A[15]), .A2(B[14]), .B1(B[15]), .B2(A[14]), .ZN(n_117));
   NOR2_X1 i_156 (.A1(n_116), .A2(n_117), .ZN(n_118));
   XNOR2_X1 i_157 (.A(n_114), .B(n_118), .ZN(n_75));
   NAND2_X1 i_158 (.A1(B[2]), .A2(A[1]), .ZN(n_119));
   NAND2_X1 i_159 (.A1(B[3]), .A2(A[2]), .ZN(n_120));
   NOR2_X1 i_160 (.A1(n_119), .A2(n_120), .ZN(n_121));
   AOI22_X1 i_161 (.A1(B[2]), .A2(A[2]), .B1(B[3]), .B2(A[1]), .ZN(n_122));
   NOR2_X1 i_162 (.A1(n_121), .A2(n_122), .ZN(n_123));
   NAND2_X1 i_163 (.A1(B[4]), .A2(A[0]), .ZN(n_124));
   XNOR2_X1 i_164 (.A(n_123), .B(n_124), .ZN(n_271));
   AND2_X1 i_165 (.A1(A[0]), .A2(B[0]), .ZN(Z[0]));
   INV_X1 i_166 (.A(n_119), .ZN(n_125));
   NAND3_X1 i_167 (.A1(n_125), .A2(B[1]), .A3(A[0]), .ZN(n_126));
   INV_X1 i_168 (.A(n_126), .ZN(n_127));
   AOI22_X1 i_169 (.A1(B[1]), .A2(A[1]), .B1(B[2]), .B2(A[0]), .ZN(n_128));
   NOR2_X1 i_170 (.A1(n_127), .A2(n_128), .ZN(n_129));
   AOI21_X1 i_171 (.A(n_129), .B1(A[2]), .B2(B[0]), .ZN(n_130));
   NAND3_X1 i_172 (.A1(Z[0]), .A2(B[1]), .A3(A[1]), .ZN(n_131));
   NAND3_X1 i_173 (.A1(n_129), .A2(A[2]), .A3(B[0]), .ZN(n_132));
   AOI21_X1 i_174 (.A(n_130), .B1(n_131), .B2(n_132), .ZN(n_76));
   NAND3_X1 i_175 (.A1(n_125), .A2(A[2]), .A3(B[1]), .ZN(n_133));
   AOI21_X1 i_176 (.A(n_125), .B1(A[2]), .B2(B[1]), .ZN(n_134));
   INV_X1 i_177 (.A(n_134), .ZN(n_135));
   NAND2_X1 i_178 (.A1(n_133), .A2(n_135), .ZN(n_136));
   NAND2_X1 i_179 (.A1(B[3]), .A2(A[0]), .ZN(n_137));
   XOR2_X1 i_180 (.A(n_136), .B(n_137), .Z(n_261));
   NAND2_X1 i_181 (.A1(A[3]), .A2(B[0]), .ZN(n_138));
   XOR2_X1 i_182 (.A(n_126), .B(n_138), .Z(n_266));
   AOI22_X1 i_183 (.A1(A[15]), .A2(B[11]), .B1(A[14]), .B2(B[12]), .ZN(n_139));
   NAND2_X1 i_184 (.A1(A[14]), .A2(B[11]), .ZN(n_140));
   INV_X1 i_185 (.A(A[15]), .ZN(n_141));
   INV_X1 i_186 (.A(B[10]), .ZN(n_142));
   OR3_X1 i_187 (.A1(n_140), .A2(n_141), .A3(n_142), .ZN(n_143));
   INV_X1 i_188 (.A(n_143), .ZN(n_144));
   AND2_X1 i_189 (.A1(A[13]), .A2(B[12]), .ZN(n_145));
   OAI21_X1 i_190 (.A(n_140), .B1(n_141), .B2(n_142), .ZN(n_146));
   AOI21_X1 i_191 (.A(n_144), .B1(n_145), .B2(n_146), .ZN(n_147));
   NAND2_X1 i_192 (.A1(A[15]), .A2(B[12]), .ZN(n_148));
   NOR2_X1 i_193 (.A1(n_140), .A2(n_148), .ZN(n_149));
   INV_X1 i_194 (.A(n_149), .ZN(n_150));
   AOI21_X1 i_195 (.A(n_139), .B1(n_147), .B2(n_150), .ZN(n_151));
   AND2_X1 i_196 (.A1(B[13]), .A2(A[12]), .ZN(n_152));
   NAND3_X1 i_197 (.A1(n_152), .A2(B[14]), .A3(A[13]), .ZN(n_153));
   AOI22_X1 i_198 (.A1(B[14]), .A2(A[12]), .B1(A[13]), .B2(B[13]), .ZN(n_154));
   NAND2_X1 i_199 (.A1(B[15]), .A2(A[11]), .ZN(n_155));
   OAI21_X1 i_200 (.A(n_153), .B1(n_154), .B2(n_155), .ZN(n_156));
   NOR2_X1 i_201 (.A1(n_151), .A2(n_156), .ZN(n_157));
   NAND2_X1 i_202 (.A1(n_151), .A2(n_156), .ZN(n_158));
   AOI21_X1 i_203 (.A(n_157), .B1(n_148), .B2(n_158), .ZN(n_77));
   NAND2_X1 i_204 (.A1(n_108), .A2(n_112), .ZN(n_159));
   XNOR2_X1 i_205 (.A(n_159), .B(n_113), .ZN(n_78));
   NAND3_X1 i_206 (.A1(n_107), .A2(A[13]), .A3(B[13]), .ZN(n_160));
   AOI22_X1 i_207 (.A1(B[14]), .A2(A[13]), .B1(A[14]), .B2(B[13]), .ZN(n_161));
   NAND2_X1 i_208 (.A1(B[15]), .A2(A[12]), .ZN(n_162));
   OAI21_X1 i_209 (.A(n_160), .B1(n_161), .B2(n_162), .ZN(n_79));
   INV_X1 i_210 (.A(n_157), .ZN(n_163));
   NAND2_X1 i_211 (.A1(n_163), .A2(n_158), .ZN(n_164));
   XOR2_X1 i_212 (.A(n_164), .B(n_148), .Z(n_80));
   INV_X1 i_213 (.A(n_161), .ZN(n_165));
   NAND2_X1 i_214 (.A1(n_160), .A2(n_165), .ZN(n_166));
   XOR2_X1 i_215 (.A(n_166), .B(n_162), .Z(n_81));
   INV_X1 i_216 (.A(n_154), .ZN(n_167));
   NAND2_X1 i_217 (.A1(n_153), .A2(n_167), .ZN(n_168));
   XOR2_X1 i_218 (.A(n_168), .B(n_155), .Z(n_82));
   NOR2_X1 i_219 (.A1(n_149), .A2(n_139), .ZN(n_169));
   XNOR2_X1 i_220 (.A(n_147), .B(n_169), .ZN(n_83));
   NAND3_X1 i_221 (.A1(n_152), .A2(B[14]), .A3(A[11]), .ZN(n_170));
   AOI21_X1 i_222 (.A(n_152), .B1(B[14]), .B2(A[11]), .ZN(n_171));
   NAND2_X1 i_223 (.A1(B[15]), .A2(A[10]), .ZN(n_172));
   OAI21_X1 i_224 (.A(n_170), .B1(n_171), .B2(n_172), .ZN(n_84));
   INV_X1 i_225 (.A(n_171), .ZN(n_173));
   NAND2_X1 i_226 (.A1(n_170), .A2(n_173), .ZN(n_174));
   XOR2_X1 i_227 (.A(n_174), .B(n_172), .Z(n_85));
   NAND2_X1 i_228 (.A1(n_143), .A2(n_146), .ZN(n_175));
   XNOR2_X1 i_229 (.A(n_175), .B(n_145), .ZN(n_86));
   NAND2_X1 i_230 (.A1(A[13]), .A2(B[10]), .ZN(n_176));
   INV_X1 i_231 (.A(n_176), .ZN(n_177));
   NAND3_X1 i_232 (.A1(n_177), .A2(A[12]), .A3(B[11]), .ZN(n_178));
   AOI21_X1 i_233 (.A(n_177), .B1(A[12]), .B2(B[11]), .ZN(n_179));
   NAND2_X1 i_234 (.A1(A[11]), .A2(B[12]), .ZN(n_180));
   OAI21_X1 i_235 (.A(n_178), .B1(n_179), .B2(n_180), .ZN(n_181));
   NAND4_X1 i_236 (.A1(B[14]), .A2(B[13]), .A3(A[10]), .A4(A[9]), .ZN(n_182));
   AOI22_X1 i_237 (.A1(B[14]), .A2(A[9]), .B1(B[13]), .B2(A[10]), .ZN(n_183));
   NAND2_X1 i_238 (.A1(B[15]), .A2(A[8]), .ZN(n_184));
   OAI21_X1 i_239 (.A(n_182), .B1(n_183), .B2(n_184), .ZN(n_185));
   NOR2_X1 i_240 (.A1(n_181), .A2(n_185), .ZN(n_186));
   NAND2_X1 i_241 (.A1(A[15]), .A2(B[9]), .ZN(n_187));
   NAND2_X1 i_242 (.A1(n_181), .A2(n_185), .ZN(n_188));
   AOI21_X1 i_243 (.A(n_186), .B1(n_187), .B2(n_188), .ZN(n_87));
   NAND4_X1 i_244 (.A1(B[14]), .A2(B[13]), .A3(A[11]), .A4(A[10]), .ZN(n_189));
   AOI22_X1 i_245 (.A1(B[14]), .A2(A[10]), .B1(B[13]), .B2(A[11]), .ZN(n_190));
   NAND2_X1 i_246 (.A1(B[15]), .A2(A[9]), .ZN(n_191));
   OAI21_X1 i_247 (.A(n_189), .B1(n_190), .B2(n_191), .ZN(n_88));
   NOR2_X1 i_248 (.A1(n_140), .A2(n_176), .ZN(n_192));
   INV_X1 i_249 (.A(n_192), .ZN(n_193));
   AOI22_X1 i_250 (.A1(A[13]), .A2(B[11]), .B1(A[14]), .B2(B[10]), .ZN(n_194));
   NAND2_X1 i_251 (.A1(A[12]), .A2(B[12]), .ZN(n_195));
   OAI21_X1 i_252 (.A(n_193), .B1(n_194), .B2(n_195), .ZN(n_89));
   INV_X1 i_253 (.A(n_186), .ZN(n_196));
   NAND2_X1 i_254 (.A1(n_188), .A2(n_196), .ZN(n_197));
   XOR2_X1 i_255 (.A(n_197), .B(n_187), .Z(n_90));
   INV_X1 i_256 (.A(n_190), .ZN(n_198));
   NAND2_X1 i_257 (.A1(n_198), .A2(n_189), .ZN(n_199));
   XOR2_X1 i_258 (.A(n_199), .B(n_191), .Z(n_91));
   NOR2_X1 i_259 (.A1(n_192), .A2(n_194), .ZN(n_200));
   XNOR2_X1 i_260 (.A(n_200), .B(n_195), .ZN(n_92));
   INV_X1 i_261 (.A(B[9]), .ZN(n_201));
   NAND2_X1 i_262 (.A1(A[14]), .A2(B[8]), .ZN(n_202));
   NAND2_X1 i_263 (.A1(A[15]), .A2(B[7]), .ZN(n_203));
   AOI211_X1 i_264 (.A(n_111), .B(n_201), .C1(n_202), .C2(n_203), .ZN(n_204));
   AOI21_X1 i_265 (.A(n_204), .B1(A[15]), .B2(B[8]), .ZN(n_205));
   INV_X1 i_266 (.A(A[14]), .ZN(n_206));
   INV_X1 i_267 (.A(B[7]), .ZN(n_207));
   NOR2_X1 i_268 (.A1(n_206), .A2(n_207), .ZN(n_208));
   OAI211_X1 i_269 (.A(A[15]), .B(B[8]), .C1(n_204), .C2(n_208), .ZN(n_209));
   NAND2_X1 i_270 (.A1(A[14]), .A2(B[9]), .ZN(n_210));
   AOI21_X1 i_271 (.A(n_205), .B1(n_209), .B2(n_210), .ZN(n_93));
   INV_X1 i_272 (.A(n_183), .ZN(n_211));
   NAND2_X1 i_273 (.A1(n_211), .A2(n_182), .ZN(n_212));
   XOR2_X1 i_274 (.A(n_212), .B(n_184), .Z(n_94));
   INV_X1 i_275 (.A(n_179), .ZN(n_213));
   NAND2_X1 i_276 (.A1(n_178), .A2(n_213), .ZN(n_214));
   XOR2_X1 i_277 (.A(n_214), .B(n_180), .Z(n_95));
   INV_X1 i_278 (.A(n_205), .ZN(n_215));
   NAND2_X1 i_279 (.A1(n_209), .A2(n_215), .ZN(n_216));
   XOR2_X1 i_280 (.A(n_216), .B(n_210), .Z(n_96));
   NAND4_X1 i_281 (.A1(B[14]), .A2(B[13]), .A3(A[8]), .A4(A[9]), .ZN(n_217));
   AOI22_X1 i_282 (.A1(B[14]), .A2(A[8]), .B1(B[13]), .B2(A[9]), .ZN(n_218));
   NAND2_X1 i_283 (.A1(B[15]), .A2(A[7]), .ZN(n_219));
   OAI21_X1 i_284 (.A(n_217), .B1(n_218), .B2(n_219), .ZN(n_97));
   NAND4_X1 i_285 (.A1(A[11]), .A2(A[12]), .A3(B[11]), .A4(B[10]), .ZN(n_220));
   AOI22_X1 i_286 (.A1(A[11]), .A2(B[11]), .B1(A[12]), .B2(B[10]), .ZN(n_221));
   NAND2_X1 i_287 (.A1(B[12]), .A2(A[10]), .ZN(n_222));
   OAI21_X1 i_288 (.A(n_220), .B1(n_221), .B2(n_222), .ZN(n_98));
   INV_X1 i_289 (.A(n_218), .ZN(n_223));
   NAND2_X1 i_290 (.A1(n_223), .A2(n_217), .ZN(n_224));
   XOR2_X1 i_291 (.A(n_224), .B(n_219), .Z(n_99));
   INV_X1 i_292 (.A(n_221), .ZN(n_225));
   NAND2_X1 i_293 (.A1(n_225), .A2(n_220), .ZN(n_226));
   XOR2_X1 i_294 (.A(n_226), .B(n_222), .Z(n_100));
   XOR2_X1 i_295 (.A(n_202), .B(n_203), .Z(n_227));
   NAND2_X1 i_296 (.A1(A[13]), .A2(B[9]), .ZN(n_228));
   XNOR2_X1 i_297 (.A(n_227), .B(n_228), .ZN(n_101));
   NAND4_X1 i_298 (.A1(B[11]), .A2(A[10]), .A3(B[10]), .A4(A[9]), .ZN(n_229));
   AOI22_X1 i_299 (.A1(B[11]), .A2(A[9]), .B1(A[10]), .B2(B[10]), .ZN(n_230));
   NAND2_X1 i_300 (.A1(B[12]), .A2(A[8]), .ZN(n_231));
   OAI21_X1 i_301 (.A(n_229), .B1(n_230), .B2(n_231), .ZN(n_232));
   NAND4_X1 i_302 (.A1(A[13]), .A2(A[12]), .A3(B[8]), .A4(B[7]), .ZN(n_233));
   AOI22_X1 i_303 (.A1(A[12]), .A2(B[8]), .B1(A[13]), .B2(B[7]), .ZN(n_234));
   NAND2_X1 i_304 (.A1(A[11]), .A2(B[9]), .ZN(n_235));
   OAI21_X1 i_305 (.A(n_233), .B1(n_234), .B2(n_235), .ZN(n_236));
   NOR2_X1 i_306 (.A1(n_232), .A2(n_236), .ZN(n_237));
   NAND2_X1 i_307 (.A1(A[15]), .A2(B[6]), .ZN(n_238));
   NAND2_X1 i_308 (.A1(n_232), .A2(n_236), .ZN(n_239));
   AOI21_X1 i_309 (.A(n_237), .B1(n_238), .B2(n_239), .ZN(n_102));
   NAND4_X1 i_310 (.A1(B[14]), .A2(B[13]), .A3(A[8]), .A4(A[7]), .ZN(n_240));
   AOI22_X1 i_311 (.A1(B[14]), .A2(A[7]), .B1(B[13]), .B2(A[8]), .ZN(n_241));
   NAND2_X1 i_312 (.A1(B[15]), .A2(A[6]), .ZN(n_242));
   OAI21_X1 i_313 (.A(n_240), .B1(n_241), .B2(n_242), .ZN(n_952));
   NAND4_X1 i_314 (.A1(A[11]), .A2(B[11]), .A3(A[10]), .A4(B[10]), .ZN(n_243));
   AOI22_X1 i_315 (.A1(B[11]), .A2(A[10]), .B1(A[11]), .B2(B[10]), .ZN(n_244));
   NAND2_X1 i_316 (.A1(B[12]), .A2(A[9]), .ZN(n_245));
   OAI21_X1 i_317 (.A(n_243), .B1(n_244), .B2(n_245), .ZN(n_959));
   OR3_X1 i_318 (.A1(n_202), .A2(n_111), .A3(n_207), .ZN(n_246));
   AOI21_X1 i_319 (.A(n_208), .B1(A[13]), .B2(B[8]), .ZN(n_247));
   NAND2_X1 i_320 (.A1(A[12]), .A2(B[9]), .ZN(n_248));
   OAI21_X1 i_321 (.A(n_246), .B1(n_247), .B2(n_248), .ZN(n_103));
   INV_X1 i_322 (.A(n_237), .ZN(n_249));
   NAND2_X1 i_323 (.A1(n_249), .A2(n_239), .ZN(n_250));
   XOR2_X1 i_324 (.A(n_250), .B(n_238), .Z(n_104));
   INV_X1 i_325 (.A(n_241), .ZN(n_251));
   NAND2_X1 i_326 (.A1(n_251), .A2(n_240), .ZN(n_252));
   XOR2_X1 i_327 (.A(n_252), .B(n_242), .Z(n_951));
   INV_X1 i_328 (.A(n_244), .ZN(n_253));
   NAND2_X1 i_329 (.A1(n_253), .A2(n_243), .ZN(n_254));
   XOR2_X1 i_330 (.A(n_254), .B(n_245), .Z(n_958));
   INV_X1 i_331 (.A(n_247), .ZN(n_255));
   NAND2_X1 i_332 (.A1(n_246), .A2(n_255), .ZN(n_256));
   XOR2_X1 i_333 (.A(n_256), .B(n_248), .Z(n_105));
   NAND4_X1 i_334 (.A1(B[14]), .A2(B[13]), .A3(A[7]), .A4(A[6]), .ZN(n_257));
   AOI22_X1 i_335 (.A1(B[14]), .A2(A[6]), .B1(B[13]), .B2(A[7]), .ZN(n_258));
   NAND2_X1 i_336 (.A1(B[15]), .A2(A[5]), .ZN(n_259));
   OAI21_X1 i_337 (.A(n_257), .B1(n_258), .B2(n_259), .ZN(n_911));
   INV_X1 i_338 (.A(n_258), .ZN(n_260));
   NAND2_X1 i_339 (.A1(n_260), .A2(n_257), .ZN(n_263));
   XOR2_X1 i_340 (.A(n_263), .B(n_259), .Z(n_910));
   INV_X1 i_341 (.A(n_230), .ZN(n_264));
   NAND2_X1 i_342 (.A1(n_264), .A2(n_229), .ZN(n_265));
   XOR2_X1 i_343 (.A(n_265), .B(n_231), .Z(n_917));
   INV_X1 i_344 (.A(n_234), .ZN(n_267));
   NAND2_X1 i_345 (.A1(n_267), .A2(n_233), .ZN(n_268));
   XOR2_X1 i_346 (.A(n_268), .B(n_235), .Z(n_924));
   INV_X1 i_347 (.A(B[6]), .ZN(n_269));
   NAND2_X1 i_348 (.A1(A[14]), .A2(B[5]), .ZN(n_270));
   NAND2_X1 i_349 (.A1(A[15]), .A2(B[4]), .ZN(n_273));
   AOI211_X1 i_350 (.A(n_111), .B(n_269), .C1(n_270), .C2(n_273), .ZN(n_274));
   INV_X1 i_351 (.A(B[4]), .ZN(n_275));
   NOR2_X1 i_352 (.A1(n_206), .A2(n_275), .ZN(n_276));
   OAI211_X1 i_353 (.A(A[15]), .B(B[5]), .C1(n_274), .C2(n_276), .ZN(n_279));
   AOI21_X1 i_354 (.A(n_274), .B1(A[15]), .B2(B[5]), .ZN(n_280));
   NAND2_X1 i_355 (.A1(A[14]), .A2(B[6]), .ZN(n_281));
   OAI21_X1 i_356 (.A(n_279), .B1(n_280), .B2(n_281), .ZN(n_931));
   AND2_X1 i_357 (.A1(n_280), .A2(n_281), .ZN(n_282));
   OAI22_X1 i_358 (.A1(n_279), .A2(n_281), .B1(n_931), .B2(n_282), .ZN(n_930));
   NAND4_X1 i_359 (.A1(B[14]), .A2(B[13]), .A3(A[5]), .A4(A[6]), .ZN(n_283));
   AOI22_X1 i_360 (.A1(B[14]), .A2(A[5]), .B1(B[13]), .B2(A[6]), .ZN(n_286));
   NAND2_X1 i_361 (.A1(B[15]), .A2(A[4]), .ZN(n_287));
   OAI21_X1 i_362 (.A(n_283), .B1(n_286), .B2(n_287), .ZN(n_869));
   NAND4_X1 i_363 (.A1(B[11]), .A2(B[10]), .A3(A[8]), .A4(A[9]), .ZN(n_289));
   AOI22_X1 i_364 (.A1(B[11]), .A2(A[8]), .B1(B[10]), .B2(A[9]), .ZN(n_290));
   NAND2_X1 i_365 (.A1(B[12]), .A2(A[7]), .ZN(n_291));
   OAI21_X1 i_366 (.A(n_289), .B1(n_290), .B2(n_291), .ZN(n_876));
   NAND4_X1 i_367 (.A1(A[11]), .A2(A[12]), .A3(B[8]), .A4(B[7]), .ZN(n_292));
   AOI22_X1 i_368 (.A1(A[11]), .A2(B[8]), .B1(A[12]), .B2(B[7]), .ZN(n_293));
   NAND2_X1 i_369 (.A1(A[10]), .A2(B[9]), .ZN(n_294));
   OAI21_X1 i_370 (.A(n_292), .B1(n_293), .B2(n_294), .ZN(n_883));
   INV_X1 i_371 (.A(n_286), .ZN(n_296));
   NAND2_X1 i_372 (.A1(n_296), .A2(n_283), .ZN(n_297));
   XOR2_X1 i_373 (.A(n_297), .B(n_287), .Z(n_868));
   INV_X1 i_374 (.A(n_290), .ZN(n_298));
   NAND2_X1 i_375 (.A1(n_298), .A2(n_289), .ZN(n_299));
   XOR2_X1 i_376 (.A(n_299), .B(n_291), .Z(n_875));
   INV_X1 i_377 (.A(n_293), .ZN(n_304));
   NAND2_X1 i_378 (.A1(n_304), .A2(n_292), .ZN(n_305));
   XOR2_X1 i_379 (.A(n_305), .B(n_294), .Z(n_882));
   XOR2_X1 i_380 (.A(n_270), .B(n_273), .Z(n_308));
   NAND2_X1 i_381 (.A1(A[13]), .A2(B[6]), .ZN(n_309));
   XNOR2_X1 i_382 (.A(n_308), .B(n_309), .ZN(n_889));
   NAND2_X1 i_383 (.A1(A[9]), .A2(B[8]), .ZN(n_310));
   INV_X1 i_384 (.A(A[10]), .ZN(n_311));
   OR3_X1 i_385 (.A1(n_310), .A2(n_311), .A3(n_207), .ZN(n_312));
   INV_X1 i_386 (.A(n_312), .ZN(n_314));
   AND2_X1 i_387 (.A1(A[8]), .A2(B[9]), .ZN(n_315));
   OAI21_X1 i_388 (.A(n_310), .B1(n_311), .B2(n_207), .ZN(n_316));
   AOI21_X1 i_389 (.A(n_314), .B1(n_315), .B2(n_316), .ZN(n_317));
   NAND2_X1 i_390 (.A1(A[12]), .A2(B[5]), .ZN(n_318));
   NAND2_X1 i_391 (.A1(A[13]), .A2(B[4]), .ZN(n_319));
   NOR2_X1 i_392 (.A1(n_318), .A2(n_319), .ZN(n_322));
   AND2_X1 i_393 (.A1(A[11]), .A2(B[6]), .ZN(n_323));
   NAND2_X1 i_394 (.A1(n_318), .A2(n_319), .ZN(n_324));
   AOI21_X1 i_395 (.A(n_322), .B1(n_323), .B2(n_324), .ZN(n_325));
   NAND2_X1 i_396 (.A1(n_317), .A2(n_325), .ZN(n_330));
   INV_X1 i_397 (.A(n_330), .ZN(n_331));
   NAND2_X1 i_398 (.A1(A[15]), .A2(B[3]), .ZN(n_334));
   OR2_X1 i_399 (.A1(n_317), .A2(n_325), .ZN(n_335));
   AOI21_X1 i_400 (.A(n_331), .B1(n_334), .B2(n_335), .ZN(n_847));
   NAND4_X1 i_401 (.A1(B[14]), .A2(B[13]), .A3(A[5]), .A4(A[4]), .ZN(n_336));
   AOI22_X1 i_402 (.A1(B[14]), .A2(A[4]), .B1(B[13]), .B2(A[5]), .ZN(n_337));
   NAND2_X1 i_403 (.A1(B[15]), .A2(A[3]), .ZN(n_338));
   OAI21_X1 i_404 (.A(n_336), .B1(n_337), .B2(n_338), .ZN(n_819));
   NAND4_X1 i_405 (.A1(B[11]), .A2(B[10]), .A3(A[8]), .A4(A[7]), .ZN(n_341));
   AOI22_X1 i_406 (.A1(B[11]), .A2(A[7]), .B1(B[10]), .B2(A[8]), .ZN(n_342));
   NAND2_X1 i_407 (.A1(B[12]), .A2(A[6]), .ZN(n_343));
   OAI21_X1 i_408 (.A(n_341), .B1(n_342), .B2(n_343), .ZN(n_826));
   NAND4_X1 i_409 (.A1(A[11]), .A2(A[10]), .A3(B[8]), .A4(B[7]), .ZN(n_344));
   AOI22_X1 i_410 (.A1(A[10]), .A2(B[8]), .B1(A[11]), .B2(B[7]), .ZN(n_347));
   NAND2_X1 i_411 (.A1(A[9]), .A2(B[9]), .ZN(n_348));
   OAI21_X1 i_412 (.A(n_344), .B1(n_347), .B2(n_348), .ZN(n_833));
   OR2_X1 i_413 (.A1(n_270), .A2(n_319), .ZN(n_349));
   AOI21_X1 i_414 (.A(n_276), .B1(A[13]), .B2(B[5]), .ZN(n_350));
   NAND2_X1 i_415 (.A1(A[12]), .A2(B[6]), .ZN(n_351));
   OAI21_X1 i_416 (.A(n_349), .B1(n_350), .B2(n_351), .ZN(n_840));
   NAND2_X1 i_417 (.A1(n_335), .A2(n_330), .ZN(n_358));
   XOR2_X1 i_418 (.A(n_358), .B(n_334), .Z(n_846));
   INV_X1 i_419 (.A(n_337), .ZN(n_359));
   NAND2_X1 i_420 (.A1(n_359), .A2(n_336), .ZN(n_362));
   XOR2_X1 i_421 (.A(n_362), .B(n_338), .Z(n_818));
   INV_X1 i_422 (.A(n_342), .ZN(n_363));
   NAND2_X1 i_423 (.A1(n_363), .A2(n_341), .ZN(n_364));
   XOR2_X1 i_424 (.A(n_364), .B(n_343), .Z(n_825));
   INV_X1 i_425 (.A(n_347), .ZN(n_365));
   NAND2_X1 i_426 (.A1(n_365), .A2(n_344), .ZN(n_366));
   XOR2_X1 i_427 (.A(n_366), .B(n_348), .Z(n_832));
   INV_X1 i_428 (.A(n_350), .ZN(n_368));
   NAND2_X1 i_429 (.A1(n_349), .A2(n_368), .ZN(n_369));
   XOR2_X1 i_430 (.A(n_369), .B(n_351), .Z(n_839));
   INV_X1 i_431 (.A(B[3]), .ZN(n_370));
   NAND2_X1 i_432 (.A1(A[14]), .A2(B[2]), .ZN(n_371));
   NAND2_X1 i_433 (.A1(A[15]), .A2(B[1]), .ZN(n_372));
   AOI211_X1 i_434 (.A(n_111), .B(n_370), .C1(n_371), .C2(n_372), .ZN(n_373));
   AOI21_X1 i_435 (.A(n_373), .B1(A[15]), .B2(B[2]), .ZN(n_375));
   AND2_X1 i_436 (.A1(A[14]), .A2(B[1]), .ZN(n_376));
   OAI211_X1 i_437 (.A(A[15]), .B(B[2]), .C1(n_373), .C2(n_376), .ZN(n_377));
   NAND2_X1 i_438 (.A1(A[14]), .A2(B[3]), .ZN(n_378));
   AOI21_X1 i_439 (.A(n_375), .B1(n_377), .B2(n_378), .ZN(n_794));
   NAND2_X1 i_440 (.A1(B[14]), .A2(A[3]), .ZN(n_387));
   INV_X1 i_441 (.A(n_387), .ZN(n_388));
   NAND3_X1 i_442 (.A1(n_388), .A2(B[13]), .A3(A[4]), .ZN(n_391));
   AOI21_X1 i_443 (.A(n_388), .B1(B[13]), .B2(A[4]), .ZN(n_392));
   NAND2_X1 i_444 (.A1(B[15]), .A2(A[2]), .ZN(n_393));
   OAI21_X1 i_445 (.A(n_391), .B1(n_392), .B2(n_393), .ZN(n_767));
   NAND2_X1 i_446 (.A1(B[11]), .A2(A[6]), .ZN(n_394));
   INV_X1 i_447 (.A(n_394), .ZN(n_395));
   NAND3_X1 i_448 (.A1(n_395), .A2(B[10]), .A3(A[7]), .ZN(n_398));
   AOI21_X1 i_449 (.A(n_395), .B1(B[10]), .B2(A[7]), .ZN(n_399));
   NAND2_X1 i_450 (.A1(B[12]), .A2(A[5]), .ZN(n_400));
   OAI21_X1 i_451 (.A(n_398), .B1(n_399), .B2(n_400), .ZN(n_774));
   INV_X1 i_452 (.A(n_392), .ZN(n_401));
   NAND2_X1 i_453 (.A1(n_391), .A2(n_401), .ZN(n_402));
   XOR2_X1 i_454 (.A(n_402), .B(n_393), .Z(n_766));
   INV_X1 i_455 (.A(n_399), .ZN(n_404));
   NAND2_X1 i_456 (.A1(n_398), .A2(n_404), .ZN(n_405));
   XOR2_X1 i_457 (.A(n_405), .B(n_400), .Z(n_773));
   NAND2_X1 i_458 (.A1(n_312), .A2(n_316), .ZN(n_406));
   XNOR2_X1 i_459 (.A(n_406), .B(n_315), .ZN(n_780));
   INV_X1 i_460 (.A(n_322), .ZN(n_407));
   NAND2_X1 i_461 (.A1(n_407), .A2(n_324), .ZN(n_408));
   XNOR2_X1 i_462 (.A(n_408), .B(n_323), .ZN(n_787));
   INV_X1 i_463 (.A(n_375), .ZN(n_409));
   NAND2_X1 i_464 (.A1(n_377), .A2(n_409), .ZN(n_412));
   XOR2_X1 i_465 (.A(n_412), .B(n_378), .Z(n_793));
   NAND2_X1 i_466 (.A1(B[13]), .A2(A[2]), .ZN(n_413));
   NOR2_X1 i_467 (.A1(n_387), .A2(n_413), .ZN(n_414));
   INV_X1 i_468 (.A(n_414), .ZN(n_415));
   AOI22_X1 i_469 (.A1(B[14]), .A2(A[2]), .B1(B[13]), .B2(A[3]), .ZN(n_424));
   NAND2_X1 i_470 (.A1(B[15]), .A2(A[1]), .ZN(n_425));
   OAI21_X1 i_471 (.A(n_415), .B1(n_424), .B2(n_425), .ZN(n_714));
   NAND2_X1 i_472 (.A1(B[10]), .A2(A[5]), .ZN(n_428));
   NOR2_X1 i_473 (.A1(n_394), .A2(n_428), .ZN(n_429));
   INV_X1 i_474 (.A(n_429), .ZN(n_430));
   AOI22_X1 i_475 (.A1(B[11]), .A2(A[5]), .B1(B[10]), .B2(A[6]), .ZN(n_431));
   NAND2_X1 i_476 (.A1(B[12]), .A2(A[4]), .ZN(n_432));
   OAI21_X1 i_477 (.A(n_430), .B1(n_431), .B2(n_432), .ZN(n_721));
   NAND2_X1 i_478 (.A1(A[8]), .A2(B[7]), .ZN(n_435));
   NOR2_X1 i_479 (.A1(n_310), .A2(n_435), .ZN(n_436));
   INV_X1 i_480 (.A(n_436), .ZN(n_437));
   AOI22_X1 i_481 (.A1(A[8]), .A2(B[8]), .B1(A[9]), .B2(B[7]), .ZN(n_438));
   NAND2_X1 i_482 (.A1(B[9]), .A2(A[7]), .ZN(n_439));
   OAI21_X1 i_483 (.A(n_437), .B1(n_438), .B2(n_439), .ZN(n_728));
   NAND2_X1 i_484 (.A1(A[11]), .A2(B[4]), .ZN(n_442));
   NOR2_X1 i_485 (.A1(n_318), .A2(n_442), .ZN(n_443));
   INV_X1 i_486 (.A(n_443), .ZN(n_444));
   AOI22_X1 i_487 (.A1(A[11]), .A2(B[5]), .B1(A[12]), .B2(B[4]), .ZN(n_445));
   NAND2_X1 i_488 (.A1(A[10]), .A2(B[6]), .ZN(n_448));
   OAI21_X1 i_489 (.A(n_444), .B1(n_445), .B2(n_448), .ZN(n_735));
   NOR2_X1 i_490 (.A1(n_414), .A2(n_424), .ZN(n_449));
   XNOR2_X1 i_491 (.A(n_449), .B(n_425), .ZN(n_713));
   NOR2_X1 i_492 (.A1(n_429), .A2(n_431), .ZN(n_450));
   XNOR2_X1 i_493 (.A(n_450), .B(n_432), .ZN(n_720));
   NOR2_X1 i_494 (.A1(n_436), .A2(n_438), .ZN(n_451));
   XNOR2_X1 i_495 (.A(n_451), .B(n_439), .ZN(n_727));
   NOR2_X1 i_496 (.A1(n_443), .A2(n_445), .ZN(n_452));
   XNOR2_X1 i_497 (.A(n_452), .B(n_448), .ZN(n_734));
   XOR2_X1 i_498 (.A(n_371), .B(n_372), .Z(n_463));
   NAND2_X1 i_499 (.A1(A[13]), .A2(B[3]), .ZN(n_464));
   XNOR2_X1 i_500 (.A(n_463), .B(n_464), .ZN(n_741));
   NAND2_X1 i_501 (.A1(A[13]), .A2(B[1]), .ZN(n_467));
   INV_X1 i_502 (.A(B[0]), .ZN(n_468));
   OR3_X1 i_503 (.A1(n_467), .A2(n_206), .A3(n_468), .ZN(n_469));
   INV_X1 i_504 (.A(n_469), .ZN(n_470));
   AND2_X1 i_505 (.A1(A[12]), .A2(B[2]), .ZN(n_471));
   OAI21_X1 i_506 (.A(n_467), .B1(n_206), .B2(n_468), .ZN(n_474));
   AOI21_X1 i_507 (.A(n_470), .B1(n_471), .B2(n_474), .ZN(n_475));
   INV_X1 i_508 (.A(n_475), .ZN(n_476));
   NAND2_X1 i_509 (.A1(A[10]), .A2(B[3]), .ZN(n_477));
   NOR2_X1 i_510 (.A1(n_442), .A2(n_477), .ZN(n_478));
   INV_X1 i_511 (.A(n_478), .ZN(n_480));
   AOI22_X1 i_512 (.A1(A[11]), .A2(B[3]), .B1(A[10]), .B2(B[4]), .ZN(n_481));
   NAND2_X1 i_513 (.A1(A[9]), .A2(B[5]), .ZN(n_482));
   OAI21_X1 i_514 (.A(n_480), .B1(n_481), .B2(n_482), .ZN(n_483));
   OR2_X1 i_515 (.A1(n_476), .A2(n_483), .ZN(n_484));
   INV_X1 i_516 (.A(n_484), .ZN(n_485));
   NAND2_X1 i_517 (.A1(A[15]), .A2(B[0]), .ZN(n_487));
   NAND2_X1 i_518 (.A1(n_476), .A2(n_483), .ZN(n_488));
   AOI21_X1 i_519 (.A(n_485), .B1(n_487), .B2(n_488), .ZN(n_690));
   INV_X1 i_520 (.A(n_413), .ZN(n_489));
   NAND3_X1 i_521 (.A1(n_489), .A2(B[14]), .A3(A[1]), .ZN(n_490));
   AOI21_X1 i_522 (.A(n_489), .B1(B[14]), .B2(A[1]), .ZN(n_503));
   NAND2_X1 i_523 (.A1(B[15]), .A2(A[0]), .ZN(n_504));
   OAI21_X1 i_524 (.A(n_490), .B1(n_503), .B2(n_504), .ZN(n_655));
   INV_X1 i_525 (.A(n_428), .ZN(n_507));
   NAND3_X1 i_526 (.A1(n_507), .A2(B[11]), .A3(A[4]), .ZN(n_508));
   AOI21_X1 i_527 (.A(n_507), .B1(B[11]), .B2(A[4]), .ZN(n_509));
   NAND2_X1 i_528 (.A1(B[12]), .A2(A[3]), .ZN(n_510));
   OAI21_X1 i_529 (.A(n_508), .B1(n_509), .B2(n_510), .ZN(n_662));
   INV_X1 i_530 (.A(n_435), .ZN(n_511));
   NAND3_X1 i_531 (.A1(n_511), .A2(B[8]), .A3(A[7]), .ZN(n_514));
   AOI21_X1 i_532 (.A(n_511), .B1(B[8]), .B2(A[7]), .ZN(n_515));
   NAND2_X1 i_533 (.A1(B[9]), .A2(A[6]), .ZN(n_516));
   OAI21_X1 i_534 (.A(n_514), .B1(n_515), .B2(n_516), .ZN(n_669));
   INV_X1 i_535 (.A(n_442), .ZN(n_517));
   NAND3_X1 i_536 (.A1(n_517), .A2(A[10]), .A3(B[5]), .ZN(n_518));
   AOI21_X1 i_537 (.A(n_517), .B1(A[10]), .B2(B[5]), .ZN(n_521));
   NAND2_X1 i_538 (.A1(A[9]), .A2(B[6]), .ZN(n_522));
   OAI21_X1 i_539 (.A(n_518), .B1(n_521), .B2(n_522), .ZN(n_676));
   OR2_X1 i_540 (.A1(n_371), .A2(n_467), .ZN(n_523));
   AOI21_X1 i_541 (.A(n_376), .B1(A[13]), .B2(B[2]), .ZN(n_524));
   NAND2_X1 i_542 (.A1(A[12]), .A2(B[3]), .ZN(n_525));
   OAI21_X1 i_543 (.A(n_523), .B1(n_524), .B2(n_525), .ZN(n_683));
   NAND2_X1 i_544 (.A1(n_488), .A2(n_484), .ZN(n_527));
   XOR2_X1 i_545 (.A(n_527), .B(n_487), .Z(n_689));
   INV_X1 i_546 (.A(n_503), .ZN(n_528));
   NAND2_X1 i_547 (.A1(n_490), .A2(n_528), .ZN(n_529));
   XOR2_X1 i_548 (.A(n_529), .B(n_504), .Z(n_654));
   INV_X1 i_549 (.A(n_509), .ZN(n_530));
   NAND2_X1 i_550 (.A1(n_508), .A2(n_530), .ZN(n_531));
   XOR2_X1 i_551 (.A(n_531), .B(n_510), .Z(n_661));
   INV_X1 i_552 (.A(n_515), .ZN(n_532));
   NAND2_X1 i_553 (.A1(n_514), .A2(n_532), .ZN(n_535));
   XOR2_X1 i_554 (.A(n_535), .B(n_516), .Z(n_668));
   INV_X1 i_555 (.A(n_521), .ZN(n_536));
   NAND2_X1 i_556 (.A1(n_518), .A2(n_536), .ZN(n_537));
   XOR2_X1 i_557 (.A(n_537), .B(n_522), .Z(n_675));
   INV_X1 i_558 (.A(n_524), .ZN(n_538));
   NAND2_X1 i_559 (.A1(n_523), .A2(n_538), .ZN(n_551));
   XOR2_X1 i_560 (.A(n_551), .B(n_525), .Z(n_682));
   NAND2_X1 i_561 (.A1(B[12]), .A2(A[1]), .ZN(n_552));
   NOR2_X1 i_562 (.A1(n_413), .A2(n_552), .ZN(n_555));
   INV_X1 i_563 (.A(n_555), .ZN(n_556));
   AOI22_X1 i_564 (.A1(B[12]), .A2(A[2]), .B1(B[13]), .B2(A[1]), .ZN(n_557));
   NAND2_X1 i_565 (.A1(B[14]), .A2(A[0]), .ZN(n_558));
   OAI21_X1 i_566 (.A(n_556), .B1(n_557), .B2(n_558), .ZN(n_604));
   NAND2_X1 i_567 (.A1(B[9]), .A2(A[4]), .ZN(n_559));
   NOR2_X1 i_568 (.A1(n_428), .A2(n_559), .ZN(n_562));
   INV_X1 i_569 (.A(n_562), .ZN(n_563));
   AOI22_X1 i_570 (.A1(B[9]), .A2(A[5]), .B1(B[10]), .B2(A[4]), .ZN(n_564));
   NAND2_X1 i_571 (.A1(B[11]), .A2(A[3]), .ZN(n_565));
   OAI21_X1 i_572 (.A(n_563), .B1(n_564), .B2(n_565), .ZN(n_611));
   NAND2_X1 i_573 (.A1(A[7]), .A2(B[6]), .ZN(n_566));
   NOR2_X1 i_574 (.A1(n_435), .A2(n_566), .ZN(n_569));
   INV_X1 i_575 (.A(n_569), .ZN(n_570));
   AOI22_X1 i_576 (.A1(A[8]), .A2(B[6]), .B1(A[7]), .B2(B[7]), .ZN(n_571));
   NAND2_X1 i_577 (.A1(B[8]), .A2(A[6]), .ZN(n_572));
   OAI21_X1 i_578 (.A(n_570), .B1(n_571), .B2(n_572), .ZN(n_618));
   NOR2_X1 i_579 (.A1(n_555), .A2(n_557), .ZN(n_573));
   XNOR2_X1 i_580 (.A(n_573), .B(n_558), .ZN(n_603));
   NOR2_X1 i_581 (.A1(n_562), .A2(n_564), .ZN(n_576));
   XNOR2_X1 i_582 (.A(n_576), .B(n_565), .ZN(n_610));
   NOR2_X1 i_583 (.A1(n_569), .A2(n_571), .ZN(n_577));
   XNOR2_X1 i_584 (.A(n_577), .B(n_572), .ZN(n_617));
   NOR2_X1 i_585 (.A1(n_478), .A2(n_481), .ZN(n_578));
   XNOR2_X1 i_586 (.A(n_578), .B(n_482), .ZN(n_624));
   NAND2_X1 i_587 (.A1(n_469), .A2(n_474), .ZN(n_579));
   XNOR2_X1 i_588 (.A(n_579), .B(n_471), .ZN(n_631));
   NAND4_X1 i_589 (.A1(A[11]), .A2(A[10]), .A3(B[2]), .A4(B[1]), .ZN(n_582));
   AOI22_X1 i_590 (.A1(A[11]), .A2(B[1]), .B1(A[10]), .B2(B[2]), .ZN(n_583));
   NAND2_X1 i_591 (.A1(A[9]), .A2(B[3]), .ZN(n_584));
   OAI21_X1 i_592 (.A(n_582), .B1(n_583), .B2(n_584), .ZN(n_585));
   AOI21_X1 i_593 (.A(n_585), .B1(A[13]), .B2(B[0]), .ZN(n_586));
   NAND2_X1 i_594 (.A1(A[12]), .A2(B[1]), .ZN(n_601));
   NAND3_X1 i_595 (.A1(n_585), .A2(A[13]), .A3(B[0]), .ZN(n_602));
   AOI21_X1 i_596 (.A(n_586), .B1(n_601), .B2(n_602), .ZN(n_581));
   INV_X1 i_597 (.A(n_552), .ZN(n_605));
   NAND3_X1 i_598 (.A1(n_605), .A2(B[11]), .A3(A[2]), .ZN(n_606));
   AOI21_X1 i_599 (.A(n_605), .B1(B[11]), .B2(A[2]), .ZN(n_607));
   NAND2_X1 i_600 (.A1(B[13]), .A2(A[0]), .ZN(n_608));
   OAI21_X1 i_601 (.A(n_606), .B1(n_607), .B2(n_608), .ZN(n_554));
   INV_X1 i_602 (.A(n_559), .ZN(n_609));
   NAND3_X1 i_603 (.A1(n_609), .A2(B[8]), .A3(A[5]), .ZN(n_612));
   AOI21_X1 i_604 (.A(n_609), .B1(B[8]), .B2(A[5]), .ZN(n_613));
   NAND2_X1 i_605 (.A1(B[10]), .A2(A[3]), .ZN(n_614));
   OAI21_X1 i_606 (.A(n_612), .B1(n_613), .B2(n_614), .ZN(n_561));
   INV_X1 i_607 (.A(n_566), .ZN(n_615));
   NAND3_X1 i_608 (.A1(n_615), .A2(A[8]), .A3(B[5]), .ZN(n_616));
   AOI21_X1 i_609 (.A(n_615), .B1(A[8]), .B2(B[5]), .ZN(n_619));
   NAND2_X1 i_610 (.A1(B[7]), .A2(A[6]), .ZN(n_620));
   OAI21_X1 i_611 (.A(n_616), .B1(n_619), .B2(n_620), .ZN(n_568));
   INV_X1 i_612 (.A(n_477), .ZN(n_621));
   NAND3_X1 i_613 (.A1(n_621), .A2(A[11]), .A3(B[2]), .ZN(n_622));
   AOI21_X1 i_614 (.A(n_621), .B1(A[11]), .B2(B[2]), .ZN(n_623));
   NAND2_X1 i_615 (.A1(A[9]), .A2(B[4]), .ZN(n_625));
   OAI21_X1 i_616 (.A(n_622), .B1(n_623), .B2(n_625), .ZN(n_575));
   INV_X1 i_617 (.A(n_607), .ZN(n_626));
   NAND2_X1 i_618 (.A1(n_606), .A2(n_626), .ZN(n_627));
   XOR2_X1 i_619 (.A(n_627), .B(n_608), .Z(n_553));
   INV_X1 i_620 (.A(n_613), .ZN(n_628));
   NAND2_X1 i_621 (.A1(n_612), .A2(n_628), .ZN(n_629));
   XOR2_X1 i_622 (.A(n_629), .B(n_614), .Z(n_560));
   INV_X1 i_623 (.A(n_619), .ZN(n_630));
   NAND2_X1 i_624 (.A1(n_616), .A2(n_630), .ZN(n_632));
   XOR2_X1 i_625 (.A(n_632), .B(n_620), .Z(n_567));
   INV_X1 i_626 (.A(n_623), .ZN(n_633));
   NAND2_X1 i_627 (.A1(n_622), .A2(n_633), .ZN(n_634));
   XOR2_X1 i_628 (.A(n_634), .B(n_625), .Z(n_574));
   INV_X1 i_629 (.A(n_586), .ZN(n_635));
   NAND2_X1 i_630 (.A1(n_635), .A2(n_602), .ZN(n_652));
   XOR2_X1 i_631 (.A(n_652), .B(n_601), .Z(n_580));
   NAND4_X1 i_632 (.A1(A[8]), .A2(A[7]), .A3(B[3]), .A4(B[4]), .ZN(n_653));
   AOI22_X1 i_633 (.A1(A[8]), .A2(B[3]), .B1(A[7]), .B2(B[4]), .ZN(n_656));
   NAND2_X1 i_634 (.A1(A[6]), .A2(B[5]), .ZN(n_657));
   OAI21_X1 i_635 (.A(n_653), .B1(n_656), .B2(n_657), .ZN(n_658));
   NAND4_X1 i_636 (.A1(A[11]), .A2(A[10]), .A3(B[1]), .A4(B[0]), .ZN(n_659));
   AOI22_X1 i_637 (.A1(A[11]), .A2(B[0]), .B1(A[10]), .B2(B[1]), .ZN(n_660));
   NAND2_X1 i_638 (.A1(A[9]), .A2(B[2]), .ZN(n_663));
   OAI21_X1 i_639 (.A(n_659), .B1(n_660), .B2(n_663), .ZN(n_664));
   NOR2_X1 i_640 (.A1(n_658), .A2(n_664), .ZN(n_665));
   NAND2_X1 i_641 (.A1(A[12]), .A2(B[0]), .ZN(n_666));
   NAND2_X1 i_642 (.A1(n_658), .A2(n_664), .ZN(n_667));
   AOI21_X1 i_643 (.A(n_665), .B1(n_666), .B2(n_667), .ZN(n_534));
   NAND4_X1 i_644 (.A1(B[11]), .A2(B[10]), .A3(A[2]), .A4(A[1]), .ZN(n_670));
   AOI22_X1 i_645 (.A1(B[10]), .A2(A[2]), .B1(B[11]), .B2(A[1]), .ZN(n_671));
   NAND2_X1 i_646 (.A1(B[12]), .A2(A[0]), .ZN(n_672));
   OAI21_X1 i_647 (.A(n_670), .B1(n_671), .B2(n_672), .ZN(n_506));
   NAND4_X1 i_648 (.A1(B[8]), .A2(B[7]), .A3(A[5]), .A4(A[4]), .ZN(n_673));
   AOI22_X1 i_649 (.A1(B[7]), .A2(A[5]), .B1(B[8]), .B2(A[4]), .ZN(n_674));
   NAND2_X1 i_650 (.A1(B[9]), .A2(A[3]), .ZN(n_677));
   OAI21_X1 i_651 (.A(n_673), .B1(n_674), .B2(n_677), .ZN(n_513));
   NAND4_X1 i_652 (.A1(A[8]), .A2(A[7]), .A3(B[4]), .A4(B[5]), .ZN(n_678));
   AOI22_X1 i_653 (.A1(A[8]), .A2(B[4]), .B1(A[7]), .B2(B[5]), .ZN(n_679));
   NAND2_X1 i_654 (.A1(A[6]), .A2(B[6]), .ZN(n_680));
   OAI21_X1 i_655 (.A(n_678), .B1(n_679), .B2(n_680), .ZN(n_520));
   INV_X1 i_656 (.A(n_665), .ZN(n_681));
   NAND2_X1 i_657 (.A1(n_681), .A2(n_667), .ZN(n_684));
   XOR2_X1 i_658 (.A(n_684), .B(n_666), .Z(n_533));
   INV_X1 i_659 (.A(n_671), .ZN(n_685));
   NAND2_X1 i_660 (.A1(n_685), .A2(n_670), .ZN(n_686));
   XOR2_X1 i_661 (.A(n_686), .B(n_672), .Z(n_505));
   INV_X1 i_662 (.A(n_674), .ZN(n_687));
   NAND2_X1 i_663 (.A1(n_687), .A2(n_673), .ZN(n_688));
   XOR2_X1 i_664 (.A(n_688), .B(n_677), .Z(n_512));
   INV_X1 i_665 (.A(n_679), .ZN(n_691));
   NAND2_X1 i_666 (.A1(n_691), .A2(n_678), .ZN(n_692));
   XOR2_X1 i_667 (.A(n_692), .B(n_680), .Z(n_519));
   INV_X1 i_668 (.A(n_583), .ZN(n_693));
   NAND2_X1 i_669 (.A1(n_693), .A2(n_582), .ZN(n_694));
   XOR2_X1 i_670 (.A(n_694), .B(n_584), .Z(n_526));
   NAND4_X1 i_671 (.A1(B[10]), .A2(B[9]), .A3(A[2]), .A4(A[1]), .ZN(n_711));
   AOI22_X1 i_672 (.A1(B[9]), .A2(A[2]), .B1(B[10]), .B2(A[1]), .ZN(n_712));
   NAND2_X1 i_673 (.A1(B[11]), .A2(A[0]), .ZN(n_715));
   OAI21_X1 i_674 (.A(n_711), .B1(n_712), .B2(n_715), .ZN(n_466));
   NAND4_X1 i_675 (.A1(B[7]), .A2(A[5]), .A3(B[6]), .A4(A[4]), .ZN(n_716));
   AOI22_X1 i_676 (.A1(A[5]), .A2(B[6]), .B1(B[7]), .B2(A[4]), .ZN(n_717));
   NAND2_X1 i_677 (.A1(B[8]), .A2(A[3]), .ZN(n_718));
   OAI21_X1 i_678 (.A(n_716), .B1(n_717), .B2(n_718), .ZN(n_473));
   INV_X1 i_679 (.A(n_712), .ZN(n_719));
   NAND2_X1 i_680 (.A1(n_719), .A2(n_711), .ZN(n_722));
   XOR2_X1 i_681 (.A(n_722), .B(n_715), .Z(n_465));
   INV_X1 i_682 (.A(n_717), .ZN(n_723));
   NAND2_X1 i_683 (.A1(n_723), .A2(n_716), .ZN(n_724));
   XOR2_X1 i_684 (.A(n_724), .B(n_718), .Z(n_472));
   INV_X1 i_685 (.A(n_656), .ZN(n_725));
   NAND2_X1 i_686 (.A1(n_725), .A2(n_653), .ZN(n_726));
   XOR2_X1 i_687 (.A(n_726), .B(n_657), .Z(n_479));
   INV_X1 i_688 (.A(n_660), .ZN(n_729));
   NAND2_X1 i_689 (.A1(n_729), .A2(n_659), .ZN(n_730));
   XOR2_X1 i_690 (.A(n_730), .B(n_663), .Z(n_486));
   NAND4_X1 i_691 (.A1(A[8]), .A2(A[7]), .A3(B[2]), .A4(B[1]), .ZN(n_731));
   AOI22_X1 i_692 (.A1(A[8]), .A2(B[1]), .B1(A[7]), .B2(B[2]), .ZN(n_732));
   NAND2_X1 i_693 (.A1(B[3]), .A2(A[6]), .ZN(n_733));
   OAI21_X1 i_694 (.A(n_731), .B1(n_732), .B2(n_733), .ZN(n_736));
   AOI21_X1 i_695 (.A(n_736), .B1(A[10]), .B2(B[0]), .ZN(n_737));
   NAND2_X1 i_696 (.A1(A[9]), .A2(B[1]), .ZN(n_738));
   NAND3_X1 i_697 (.A1(n_736), .A2(A[10]), .A3(B[0]), .ZN(n_739));
   AOI21_X1 i_698 (.A(n_737), .B1(n_738), .B2(n_739), .ZN(n_447));
   NAND4_X1 i_699 (.A1(B[9]), .A2(B[8]), .A3(A[2]), .A4(A[1]), .ZN(n_740));
   AOI22_X1 i_700 (.A1(B[8]), .A2(A[2]), .B1(B[9]), .B2(A[1]), .ZN(n_742));
   NAND2_X1 i_701 (.A1(B[10]), .A2(A[0]), .ZN(n_743));
   OAI21_X1 i_702 (.A(n_740), .B1(n_742), .B2(n_743), .ZN(n_427));
   NAND4_X1 i_703 (.A1(A[5]), .A2(B[6]), .A3(B[5]), .A4(A[4]), .ZN(n_744));
   AOI22_X1 i_704 (.A1(A[5]), .A2(B[5]), .B1(B[6]), .B2(A[4]), .ZN(n_745));
   NAND2_X1 i_705 (.A1(B[7]), .A2(A[3]), .ZN(n_764));
   OAI21_X1 i_706 (.A(n_744), .B1(n_745), .B2(n_764), .ZN(n_434));
   NAND4_X1 i_707 (.A1(A[8]), .A2(A[7]), .A3(B[3]), .A4(B[2]), .ZN(n_765));
   AOI22_X1 i_708 (.A1(A[8]), .A2(B[2]), .B1(A[7]), .B2(B[3]), .ZN(n_768));
   NAND2_X1 i_709 (.A1(A[6]), .A2(B[4]), .ZN(n_769));
   OAI21_X1 i_710 (.A(n_765), .B1(n_768), .B2(n_769), .ZN(n_441));
   INV_X1 i_711 (.A(n_742), .ZN(n_770));
   NAND2_X1 i_712 (.A1(n_770), .A2(n_740), .ZN(n_771));
   XOR2_X1 i_713 (.A(n_771), .B(n_743), .Z(n_426));
   INV_X1 i_714 (.A(n_745), .ZN(n_772));
   NAND2_X1 i_715 (.A1(n_772), .A2(n_744), .ZN(n_775));
   XOR2_X1 i_716 (.A(n_775), .B(n_764), .Z(n_433));
   INV_X1 i_717 (.A(n_768), .ZN(n_776));
   NAND2_X1 i_718 (.A1(n_776), .A2(n_765), .ZN(n_777));
   XOR2_X1 i_719 (.A(n_777), .B(n_769), .Z(n_440));
   INV_X1 i_720 (.A(n_737), .ZN(n_778));
   NAND2_X1 i_721 (.A1(n_778), .A2(n_739), .ZN(n_779));
   XOR2_X1 i_722 (.A(n_779), .B(n_738), .Z(n_446));
   NAND4_X1 i_723 (.A1(B[3]), .A2(A[5]), .A3(B[4]), .A4(A[4]), .ZN(n_781));
   AOI22_X1 i_724 (.A1(B[3]), .A2(A[5]), .B1(B[4]), .B2(A[4]), .ZN(n_782));
   NAND2_X1 i_725 (.A1(B[5]), .A2(A[3]), .ZN(n_783));
   OAI21_X1 i_726 (.A(n_781), .B1(n_782), .B2(n_783), .ZN(n_784));
   NAND4_X1 i_727 (.A1(A[8]), .A2(A[7]), .A3(B[1]), .A4(B[0]), .ZN(n_785));
   AOI22_X1 i_728 (.A1(A[8]), .A2(B[0]), .B1(A[7]), .B2(B[1]), .ZN(n_786));
   NAND2_X1 i_729 (.A1(B[2]), .A2(A[6]), .ZN(n_788));
   OAI21_X1 i_730 (.A(n_785), .B1(n_786), .B2(n_788), .ZN(n_789));
   NOR2_X1 i_731 (.A1(n_784), .A2(n_789), .ZN(n_790));
   NAND2_X1 i_732 (.A1(A[9]), .A2(B[0]), .ZN(n_791));
   NAND2_X1 i_733 (.A1(n_784), .A2(n_789), .ZN(n_792));
   AOI21_X1 i_734 (.A(n_790), .B1(n_791), .B2(n_792), .ZN(n_411));
   NAND4_X1 i_735 (.A1(B[8]), .A2(B[7]), .A3(A[2]), .A4(A[1]), .ZN(n_795));
   AOI22_X1 i_736 (.A1(B[7]), .A2(A[2]), .B1(B[8]), .B2(A[1]), .ZN(n_796));
   NAND2_X1 i_737 (.A1(B[9]), .A2(A[0]), .ZN(n_797));
   OAI21_X1 i_738 (.A(n_795), .B1(n_796), .B2(n_797), .ZN(n_390));
   NAND4_X1 i_739 (.A1(A[5]), .A2(B[4]), .A3(B[5]), .A4(A[4]), .ZN(n_798));
   AOI22_X1 i_740 (.A1(A[5]), .A2(B[4]), .B1(B[5]), .B2(A[4]), .ZN(n_799));
   NAND2_X1 i_741 (.A1(B[6]), .A2(A[3]), .ZN(n_816));
   OAI21_X1 i_742 (.A(n_798), .B1(n_799), .B2(n_816), .ZN(n_397));
   INV_X1 i_743 (.A(n_790), .ZN(n_817));
   NAND2_X1 i_744 (.A1(n_817), .A2(n_792), .ZN(n_820));
   XOR2_X1 i_745 (.A(n_820), .B(n_791), .Z(n_410));
   INV_X1 i_746 (.A(n_796), .ZN(n_821));
   NAND2_X1 i_747 (.A1(n_821), .A2(n_795), .ZN(n_822));
   XOR2_X1 i_748 (.A(n_822), .B(n_797), .Z(n_389));
   INV_X1 i_749 (.A(n_799), .ZN(n_823));
   NAND2_X1 i_750 (.A1(n_823), .A2(n_798), .ZN(n_824));
   XOR2_X1 i_751 (.A(n_824), .B(n_816), .Z(n_396));
   INV_X1 i_752 (.A(n_732), .ZN(n_827));
   NAND2_X1 i_753 (.A1(n_827), .A2(n_731), .ZN(n_828));
   XOR2_X1 i_754 (.A(n_828), .B(n_733), .Z(n_403));
   NAND4_X1 i_755 (.A1(B[7]), .A2(B[6]), .A3(A[2]), .A4(A[1]), .ZN(n_829));
   AOI22_X1 i_756 (.A1(B[6]), .A2(A[2]), .B1(B[7]), .B2(A[1]), .ZN(n_830));
   NAND2_X1 i_757 (.A1(B[8]), .A2(A[0]), .ZN(n_831));
   OAI21_X1 i_758 (.A(n_829), .B1(n_830), .B2(n_831), .ZN(n_361));
   INV_X1 i_759 (.A(n_830), .ZN(n_834));
   NAND2_X1 i_760 (.A1(n_834), .A2(n_829), .ZN(n_835));
   XOR2_X1 i_761 (.A(n_835), .B(n_831), .Z(n_360));
   INV_X1 i_762 (.A(n_782), .ZN(n_836));
   NAND2_X1 i_763 (.A1(n_836), .A2(n_781), .ZN(n_837));
   XOR2_X1 i_764 (.A(n_837), .B(n_783), .Z(n_367));
   INV_X1 i_765 (.A(n_786), .ZN(n_838));
   NAND2_X1 i_766 (.A1(n_838), .A2(n_785), .ZN(n_841));
   XOR2_X1 i_767 (.A(n_841), .B(n_788), .Z(n_374));
   NAND2_X1 i_768 (.A1(A[4]), .A2(B[1]), .ZN(n_842));
   NAND2_X1 i_769 (.A1(B[2]), .A2(A[5]), .ZN(n_843));
   NOR2_X1 i_770 (.A1(n_842), .A2(n_843), .ZN(n_844));
   INV_X1 i_771 (.A(n_844), .ZN(n_845));
   AOI22_X1 i_772 (.A1(A[5]), .A2(B[1]), .B1(B[2]), .B2(A[4]), .ZN(n_848));
   NAND2_X1 i_773 (.A1(B[3]), .A2(A[3]), .ZN(n_849));
   OAI21_X1 i_774 (.A(n_845), .B1(n_848), .B2(n_849), .ZN(n_850));
   AOI21_X1 i_775 (.A(n_850), .B1(A[7]), .B2(B[0]), .ZN(n_851));
   NAND2_X1 i_776 (.A1(A[6]), .A2(B[1]), .ZN(n_866));
   NAND3_X1 i_777 (.A1(n_850), .A2(A[7]), .A3(B[0]), .ZN(n_867));
   AOI21_X1 i_778 (.A(n_851), .B1(n_866), .B2(n_867), .ZN(n_346));
   NAND4_X1 i_779 (.A1(B[6]), .A2(A[2]), .A3(B[5]), .A4(A[1]), .ZN(n_870));
   AOI22_X1 i_780 (.A1(A[2]), .A2(B[5]), .B1(B[6]), .B2(A[1]), .ZN(n_871));
   NAND2_X1 i_781 (.A1(B[7]), .A2(A[0]), .ZN(n_872));
   OAI21_X1 i_782 (.A(n_870), .B1(n_871), .B2(n_872), .ZN(n_333));
   INV_X1 i_783 (.A(n_843), .ZN(n_873));
   NAND3_X1 i_784 (.A1(n_873), .A2(B[3]), .A3(A[4]), .ZN(n_874));
   AOI21_X1 i_785 (.A(n_873), .B1(B[3]), .B2(A[4]), .ZN(n_877));
   NAND2_X1 i_786 (.A1(B[4]), .A2(A[3]), .ZN(n_878));
   OAI21_X1 i_787 (.A(n_874), .B1(n_877), .B2(n_878), .ZN(n_340));
   INV_X1 i_788 (.A(n_871), .ZN(n_879));
   NAND2_X1 i_789 (.A1(n_879), .A2(n_870), .ZN(n_880));
   XOR2_X1 i_790 (.A(n_880), .B(n_872), .Z(n_332));
   INV_X1 i_791 (.A(n_877), .ZN(n_881));
   NAND2_X1 i_792 (.A1(n_874), .A2(n_881), .ZN(n_884));
   XOR2_X1 i_793 (.A(n_884), .B(n_878), .Z(n_339));
   INV_X1 i_794 (.A(n_851), .ZN(n_885));
   NAND2_X1 i_795 (.A1(n_885), .A2(n_867), .ZN(n_886));
   XOR2_X1 i_796 (.A(n_886), .B(n_866), .Z(n_345));
   INV_X1 i_797 (.A(A[1]), .ZN(n_887));
   OR3_X1 i_798 (.A1(n_120), .A2(n_275), .A3(n_887), .ZN(n_888));
   INV_X1 i_799 (.A(n_888), .ZN(n_890));
   AND2_X1 i_800 (.A1(B[5]), .A2(A[0]), .ZN(n_891));
   OAI21_X1 i_801 (.A(n_120), .B1(n_275), .B2(n_887), .ZN(n_892));
   AOI21_X1 i_802 (.A(n_890), .B1(n_891), .B2(n_892), .ZN(n_893));
   INV_X1 i_803 (.A(A[5]), .ZN(n_908));
   OR3_X1 i_804 (.A1(n_842), .A2(n_908), .A3(n_468), .ZN(n_909));
   INV_X1 i_805 (.A(n_909), .ZN(n_912));
   AND2_X1 i_806 (.A1(B[2]), .A2(A[3]), .ZN(n_913));
   OAI21_X1 i_807 (.A(n_842), .B1(n_908), .B2(n_468), .ZN(n_914));
   AOI21_X1 i_808 (.A(n_912), .B1(n_913), .B2(n_914), .ZN(n_915));
   NAND2_X1 i_809 (.A1(n_893), .A2(n_915), .ZN(n_916));
   INV_X1 i_810 (.A(n_916), .ZN(n_918));
   NAND2_X1 i_811 (.A1(A[6]), .A2(B[0]), .ZN(n_919));
   OR2_X1 i_812 (.A1(n_893), .A2(n_915), .ZN(n_920));
   AOI21_X1 i_813 (.A(n_918), .B1(n_919), .B2(n_920), .ZN(n_321));
   NAND4_X1 i_814 (.A1(B[4]), .A2(A[2]), .A3(B[5]), .A4(A[1]), .ZN(n_921));
   AOI22_X1 i_815 (.A1(B[4]), .A2(A[2]), .B1(B[5]), .B2(A[1]), .ZN(n_922));
   NAND2_X1 i_816 (.A1(B[6]), .A2(A[0]), .ZN(n_923));
   OAI21_X1 i_817 (.A(n_921), .B1(n_922), .B2(n_923), .ZN(n_307));
   NAND2_X1 i_818 (.A1(n_920), .A2(n_916), .ZN(n_925));
   XOR2_X1 i_819 (.A(n_925), .B(n_919), .Z(n_320));
   INV_X1 i_820 (.A(n_922), .ZN(n_926));
   NAND2_X1 i_821 (.A1(n_926), .A2(n_921), .ZN(n_927));
   XOR2_X1 i_822 (.A(n_927), .B(n_923), .Z(n_306));
   NOR2_X1 i_823 (.A1(n_844), .A2(n_848), .ZN(n_928));
   XNOR2_X1 i_824 (.A(n_928), .B(n_849), .ZN(n_313));
   NAND2_X1 i_825 (.A1(n_888), .A2(n_892), .ZN(n_929));
   XNOR2_X1 i_826 (.A(n_929), .B(n_891), .ZN(n_288));
   NAND2_X1 i_827 (.A1(n_909), .A2(n_914), .ZN(n_932));
   XNOR2_X1 i_828 (.A(n_932), .B(n_913), .ZN(n_295));
   INV_X1 i_829 (.A(n_121), .ZN(n_933));
   AOI21_X1 i_830 (.A(n_122), .B1(n_933), .B2(n_124), .ZN(n_272));
   AOI21_X1 i_831 (.A(n_138), .B1(n_126), .B2(n_842), .ZN(n_278));
   AOI22_X1 i_832 (.A1(A[3]), .A2(B[1]), .B1(A[4]), .B2(B[0]), .ZN(n_934));
   NAND3_X1 i_833 (.A1(A[4]), .A2(A[3]), .A3(B[0]), .ZN(n_935));
   OAI22_X1 i_834 (.A1(n_278), .A2(n_934), .B1(n_126), .B2(n_935), .ZN(n_277));
   OAI21_X1 i_835 (.A(n_133), .B1(n_134), .B2(n_137), .ZN(n_262));
   INV_X1 i_836 (.A(n_131), .ZN(n_936));
   AOI22_X1 i_837 (.A1(B[1]), .A2(A[0]), .B1(B[0]), .B2(A[1]), .ZN(n_949));
   NOR2_X1 i_838 (.A1(n_936), .A2(n_949), .ZN(Z[1]));
   INV_X1 i_839 (.A(n_130), .ZN(n_950));
   NAND2_X1 i_840 (.A1(n_950), .A2(n_132), .ZN(n_953));
   XOR2_X1 i_841 (.A(n_953), .B(n_131), .Z(Z[2]));
   INV_X1 i_842 (.A(n_116), .ZN(n_954));
   OAI21_X1 i_843 (.A(n_954), .B1(n_114), .B2(n_117), .ZN(n_955));
   INV_X1 i_844 (.A(n_115), .ZN(n_956));
   NAND2_X1 i_845 (.A1(n_956), .A2(n_74), .ZN(n_957));
   NOR2_X1 i_846 (.A1(n_956), .A2(n_74), .ZN(n_960));
   INV_X1 i_847 (.A(n_960), .ZN(n_961));
   NAND2_X1 i_848 (.A1(n_957), .A2(n_961), .ZN(n_962));
   XNOR2_X1 i_849 (.A(n_955), .B(n_962), .ZN(Z[30]));
   INV_X1 i_850 (.A(n_955), .ZN(n_963));
   OAI21_X1 i_851 (.A(n_957), .B1(n_963), .B2(n_960), .ZN(Z[31]));
endmodule

module multiplyOperator(A, B, Z);
   input [15:0]A;
   input [15:0]B;
   output [31:0]Z;

   datapath i_0_0 (.B(B), .A(A), .Z(Z));
endmodule

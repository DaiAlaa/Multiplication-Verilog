/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu May  6 02:00:04 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 4170347804 */

module multiplyShiftAdd(A, B, Z);
   input [3:0]A;
   input [3:0]B;
   output [7:0]Z;

   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;

   HA_X1 i_0_0_0 (.A(n_0_0_18), .B(n_0_0_21), .CO(n_0_0_1), .S(n_0_0_0));
   FA_X1 i_0_0_1 (.A(n_0_0_19), .B(n_0_0_22), .CI(n_0_0_25), .CO(n_0_0_3), 
      .S(n_0_0_2));
   HA_X1 i_0_0_2 (.A(n_0_0_31), .B(n_0_0_1), .CO(n_0_0_5), .S(n_0_0_4));
   FA_X1 i_0_0_3 (.A(n_0_0_20), .B(n_0_0_23), .CI(n_0_0_26), .CO(n_0_0_7), 
      .S(n_0_0_6));
   HA_X1 i_0_0_4 (.A(n_0_0_5), .B(n_0_0_3), .CO(n_0_0_9), .S(n_0_0_8));
   FA_X1 i_0_0_5 (.A(n_0_0_24), .B(n_0_0_27), .CI(n_0_0_7), .CO(n_0_0_11), 
      .S(n_0_0_10));
   HA_X1 i_0_0_6 (.A(n_0_0_17), .B(n_0_0_29), .CO(n_0_0_12), .S(Z[1]));
   FA_X1 i_0_0_7 (.A(n_0_0_30), .B(n_0_0_0), .CI(n_0_0_12), .CO(n_0_0_13), 
      .S(Z[2]));
   FA_X1 i_0_0_8 (.A(n_0_0_4), .B(n_0_0_2), .CI(n_0_0_13), .CO(n_0_0_14), 
      .S(Z[3]));
   FA_X1 i_0_0_9 (.A(n_0_0_8), .B(n_0_0_6), .CI(n_0_0_14), .CO(n_0_0_15), 
      .S(Z[4]));
   FA_X1 i_0_0_10 (.A(n_0_0_9), .B(n_0_0_10), .CI(n_0_0_15), .CO(n_0_0_16), 
      .S(Z[5]));
   FA_X1 i_0_0_11 (.A(n_0_0_28), .B(n_0_0_11), .CI(n_0_0_16), .CO(Z[7]), 
      .S(Z[6]));
   AND2_X1 i_0_0_12 (.A1(B[1]), .A2(A[0]), .ZN(n_0_0_17));
   AND2_X1 i_0_0_13 (.A1(B[1]), .A2(A[1]), .ZN(n_0_0_18));
   AND2_X1 i_0_0_14 (.A1(B[1]), .A2(A[2]), .ZN(n_0_0_19));
   AND2_X1 i_0_0_15 (.A1(B[1]), .A2(A[3]), .ZN(n_0_0_20));
   AND2_X1 i_0_0_16 (.A1(B[2]), .A2(A[0]), .ZN(n_0_0_21));
   AND2_X1 i_0_0_17 (.A1(B[2]), .A2(A[1]), .ZN(n_0_0_22));
   AND2_X1 i_0_0_18 (.A1(B[2]), .A2(A[2]), .ZN(n_0_0_23));
   AND2_X1 i_0_0_19 (.A1(B[2]), .A2(A[3]), .ZN(n_0_0_24));
   AND2_X1 i_0_0_20 (.A1(B[3]), .A2(A[0]), .ZN(n_0_0_25));
   AND2_X1 i_0_0_21 (.A1(B[3]), .A2(A[1]), .ZN(n_0_0_26));
   AND2_X1 i_0_0_22 (.A1(B[3]), .A2(A[2]), .ZN(n_0_0_27));
   AND2_X1 i_0_0_23 (.A1(B[3]), .A2(A[3]), .ZN(n_0_0_28));
   AND2_X1 i_0_0_24 (.A1(B[0]), .A2(A[0]), .ZN(Z[0]));
   AND2_X1 i_0_0_25 (.A1(B[0]), .A2(A[1]), .ZN(n_0_0_29));
   AND2_X1 i_0_0_26 (.A1(B[0]), .A2(A[2]), .ZN(n_0_0_30));
   AND2_X1 i_0_0_27 (.A1(B[0]), .A2(A[3]), .ZN(n_0_0_31));
endmodule

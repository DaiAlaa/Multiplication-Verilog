/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu May  6 02:01:20 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2647265133 */

module datapath(p_0, p_1, p_2, p_3, p_4, p_5, p_6, p_7, p_8, p_9, p_10, p_11, 
      p_12, p_13, p_14, p_15, sum_reg);
   input [31:0]p_0;
   input [31:0]p_1;
   input [31:0]p_2;
   input [31:0]p_3;
   input [31:0]p_4;
   input [31:0]p_5;
   input [31:0]p_6;
   input [31:0]p_7;
   input [31:0]p_8;
   input [31:0]p_9;
   input [31:0]p_10;
   input [31:0]p_11;
   input [31:0]p_12;
   input [31:0]p_13;
   input [31:0]p_14;
   input [31:0]p_15;
   output [31:0]sum_reg;

   HA_X1 i_0 (.A(p_0[2]), .B(p_1[2]), .CO(n_1), .S(n_0));
   FA_X1 i_1 (.A(p_0[3]), .B(p_1[3]), .CI(p_2[3]), .CO(n_3), .S(n_2));
   HA_X1 i_2 (.A(p_15[3]), .B(n_1), .CO(n_5), .S(n_4));
   FA_X1 i_3 (.A(p_0[4]), .B(p_1[4]), .CI(p_2[4]), .CO(n_7), .S(n_6));
   FA_X1 i_4 (.A(p_3[4]), .B(p_15[4]), .CI(n_5), .CO(n_9), .S(n_8));
   HA_X1 i_5 (.A(n_3), .B(n_8), .CO(n_11), .S(n_10));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(p_2[5]), .CO(n_13), .S(n_12));
   FA_X1 i_7 (.A(p_3[5]), .B(p_4[5]), .CI(p_15[5]), .CO(n_15), .S(n_14));
   FA_X1 i_8 (.A(n_7), .B(n_9), .CI(n_14), .CO(n_17), .S(n_16));
   HA_X1 i_9 (.A(n_12), .B(n_11), .CO(n_19), .S(n_18));
   FA_X1 i_10 (.A(p_0[6]), .B(p_1[6]), .CI(p_2[6]), .CO(n_21), .S(n_20));
   FA_X1 i_11 (.A(p_3[6]), .B(p_4[6]), .CI(p_5[6]), .CO(n_23), .S(n_22));
   FA_X1 i_12 (.A(p_15[6]), .B(n_15), .CI(n_13), .CO(n_25), .S(n_24));
   FA_X1 i_13 (.A(n_22), .B(n_20), .CI(n_24), .CO(n_27), .S(n_26));
   HA_X1 i_14 (.A(n_19), .B(n_17), .CO(n_29), .S(n_28));
   FA_X1 i_15 (.A(p_0[7]), .B(p_1[7]), .CI(p_2[7]), .CO(n_31), .S(n_30));
   FA_X1 i_16 (.A(p_3[7]), .B(p_4[7]), .CI(p_5[7]), .CO(n_33), .S(n_32));
   FA_X1 i_17 (.A(p_6[7]), .B(p_15[7]), .CI(n_23), .CO(n_35), .S(n_34));
   FA_X1 i_18 (.A(n_21), .B(n_25), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_19 (.A(n_32), .B(n_30), .CI(n_29), .CO(n_39), .S(n_38));
   HA_X1 i_20 (.A(n_36), .B(n_27), .CO(n_41), .S(n_40));
   FA_X1 i_21 (.A(p_0[8]), .B(p_1[8]), .CI(p_2[8]), .CO(n_43), .S(n_42));
   FA_X1 i_22 (.A(p_3[8]), .B(p_4[8]), .CI(p_5[8]), .CO(n_45), .S(n_44));
   FA_X1 i_23 (.A(p_6[8]), .B(p_7[8]), .CI(p_15[8]), .CO(n_47), .S(n_46));
   FA_X1 i_24 (.A(n_33), .B(n_31), .CI(n_35), .CO(n_49), .S(n_48));
   FA_X1 i_25 (.A(n_46), .B(n_44), .CI(n_42), .CO(n_51), .S(n_50));
   FA_X1 i_26 (.A(n_48), .B(n_37), .CI(n_41), .CO(n_53), .S(n_52));
   HA_X1 i_27 (.A(n_39), .B(n_50), .CO(n_55), .S(n_54));
   FA_X1 i_28 (.A(p_0[9]), .B(p_1[9]), .CI(p_2[9]), .CO(n_57), .S(n_56));
   FA_X1 i_29 (.A(p_3[9]), .B(p_4[9]), .CI(p_5[9]), .CO(n_59), .S(n_58));
   FA_X1 i_30 (.A(p_6[9]), .B(p_7[9]), .CI(p_8[9]), .CO(n_61), .S(n_60));
   FA_X1 i_31 (.A(p_15[9]), .B(n_47), .CI(n_45), .CO(n_63), .S(n_62));
   FA_X1 i_32 (.A(n_43), .B(n_60), .CI(n_58), .CO(n_65), .S(n_64));
   FA_X1 i_33 (.A(n_56), .B(n_49), .CI(n_62), .CO(n_67), .S(n_66));
   FA_X1 i_34 (.A(n_51), .B(n_64), .CI(n_66), .CO(n_69), .S(n_68));
   HA_X1 i_35 (.A(n_55), .B(n_53), .CO(n_71), .S(n_70));
   FA_X1 i_36 (.A(p_0[10]), .B(p_1[10]), .CI(p_2[10]), .CO(n_73), .S(n_72));
   FA_X1 i_37 (.A(p_3[10]), .B(p_4[10]), .CI(p_5[10]), .CO(n_75), .S(n_74));
   FA_X1 i_38 (.A(p_6[10]), .B(p_7[10]), .CI(p_8[10]), .CO(n_77), .S(n_76));
   FA_X1 i_39 (.A(p_9[10]), .B(p_15[10]), .CI(n_61), .CO(n_79), .S(n_78));
   FA_X1 i_40 (.A(n_59), .B(n_57), .CI(n_63), .CO(n_81), .S(n_80));
   FA_X1 i_41 (.A(n_78), .B(n_76), .CI(n_74), .CO(n_83), .S(n_82));
   FA_X1 i_42 (.A(n_72), .B(n_80), .CI(n_65), .CO(n_85), .S(n_84));
   FA_X1 i_43 (.A(n_67), .B(n_82), .CI(n_84), .CO(n_87), .S(n_86));
   HA_X1 i_44 (.A(n_71), .B(n_69), .CO(n_89), .S(n_88));
   FA_X1 i_45 (.A(p_0[11]), .B(p_1[11]), .CI(p_2[11]), .CO(n_91), .S(n_90));
   FA_X1 i_46 (.A(p_3[11]), .B(p_4[11]), .CI(p_5[11]), .CO(n_93), .S(n_92));
   FA_X1 i_47 (.A(p_6[11]), .B(p_7[11]), .CI(p_8[11]), .CO(n_95), .S(n_94));
   FA_X1 i_48 (.A(p_9[11]), .B(p_10[11]), .CI(p_15[11]), .CO(n_97), .S(n_96));
   FA_X1 i_49 (.A(n_77), .B(n_75), .CI(n_73), .CO(n_99), .S(n_98));
   FA_X1 i_50 (.A(n_79), .B(n_96), .CI(n_94), .CO(n_101), .S(n_100));
   FA_X1 i_51 (.A(n_92), .B(n_90), .CI(n_81), .CO(n_103), .S(n_102));
   FA_X1 i_52 (.A(n_98), .B(n_83), .CI(n_85), .CO(n_105), .S(n_104));
   FA_X1 i_53 (.A(n_102), .B(n_100), .CI(n_104), .CO(n_107), .S(n_106));
   HA_X1 i_54 (.A(n_89), .B(n_87), .CO(n_109), .S(n_108));
   FA_X1 i_55 (.A(p_0[12]), .B(p_1[12]), .CI(p_2[12]), .CO(n_111), .S(n_110));
   FA_X1 i_56 (.A(p_3[12]), .B(p_4[12]), .CI(p_5[12]), .CO(n_113), .S(n_112));
   FA_X1 i_57 (.A(p_6[12]), .B(p_7[12]), .CI(p_8[12]), .CO(n_115), .S(n_114));
   FA_X1 i_58 (.A(p_9[12]), .B(p_10[12]), .CI(p_11[12]), .CO(n_117), .S(n_116));
   FA_X1 i_59 (.A(p_15[12]), .B(n_97), .CI(n_95), .CO(n_119), .S(n_118));
   FA_X1 i_60 (.A(n_93), .B(n_91), .CI(n_99), .CO(n_121), .S(n_120));
   FA_X1 i_61 (.A(n_116), .B(n_114), .CI(n_112), .CO(n_123), .S(n_122));
   FA_X1 i_62 (.A(n_110), .B(n_120), .CI(n_118), .CO(n_125), .S(n_124));
   FA_X1 i_63 (.A(n_101), .B(n_103), .CI(n_122), .CO(n_127), .S(n_126));
   FA_X1 i_64 (.A(n_105), .B(n_124), .CI(n_126), .CO(n_129), .S(n_128));
   HA_X1 i_65 (.A(n_107), .B(n_109), .CO(n_131), .S(n_130));
   FA_X1 i_66 (.A(p_0[13]), .B(p_1[13]), .CI(p_2[13]), .CO(n_133), .S(n_132));
   FA_X1 i_67 (.A(p_3[13]), .B(p_4[13]), .CI(p_5[13]), .CO(n_135), .S(n_134));
   FA_X1 i_68 (.A(p_6[13]), .B(p_7[13]), .CI(p_8[13]), .CO(n_137), .S(n_136));
   FA_X1 i_69 (.A(p_9[13]), .B(p_10[13]), .CI(p_11[13]), .CO(n_139), .S(n_138));
   FA_X1 i_70 (.A(p_12[13]), .B(p_15[13]), .CI(n_117), .CO(n_141), .S(n_140));
   FA_X1 i_71 (.A(n_115), .B(n_113), .CI(n_111), .CO(n_143), .S(n_142));
   FA_X1 i_72 (.A(n_119), .B(n_140), .CI(n_138), .CO(n_145), .S(n_144));
   FA_X1 i_73 (.A(n_136), .B(n_134), .CI(n_132), .CO(n_147), .S(n_146));
   FA_X1 i_74 (.A(n_121), .B(n_142), .CI(n_123), .CO(n_149), .S(n_148));
   FA_X1 i_75 (.A(n_125), .B(n_146), .CI(n_144), .CO(n_151), .S(n_150));
   FA_X1 i_76 (.A(n_148), .B(n_127), .CI(n_129), .CO(n_153), .S(n_152));
   HA_X1 i_77 (.A(n_150), .B(n_131), .CO(n_155), .S(n_154));
   FA_X1 i_78 (.A(p_0[14]), .B(p_1[14]), .CI(p_2[14]), .CO(n_157), .S(n_156));
   FA_X1 i_79 (.A(p_3[14]), .B(p_4[14]), .CI(p_5[14]), .CO(n_159), .S(n_158));
   FA_X1 i_80 (.A(p_6[14]), .B(p_7[14]), .CI(p_8[14]), .CO(n_161), .S(n_160));
   FA_X1 i_81 (.A(p_9[14]), .B(p_10[14]), .CI(p_11[14]), .CO(n_163), .S(n_162));
   FA_X1 i_82 (.A(p_12[14]), .B(p_13[14]), .CI(p_15[14]), .CO(n_165), .S(n_164));
   FA_X1 i_83 (.A(n_139), .B(n_137), .CI(n_135), .CO(n_167), .S(n_166));
   FA_X1 i_84 (.A(n_133), .B(n_143), .CI(n_141), .CO(n_169), .S(n_168));
   FA_X1 i_85 (.A(n_164), .B(n_162), .CI(n_160), .CO(n_171), .S(n_170));
   FA_X1 i_86 (.A(n_158), .B(n_156), .CI(n_166), .CO(n_173), .S(n_172));
   FA_X1 i_87 (.A(n_147), .B(n_145), .CI(n_168), .CO(n_175), .S(n_174));
   FA_X1 i_88 (.A(n_149), .B(n_172), .CI(n_170), .CO(n_177), .S(n_176));
   FA_X1 i_89 (.A(n_174), .B(n_151), .CI(n_176), .CO(n_179), .S(n_178));
   HA_X1 i_90 (.A(n_153), .B(n_155), .CO(n_181), .S(n_180));
   FA_X1 i_91 (.A(p_0[15]), .B(p_1[15]), .CI(p_2[15]), .CO(n_183), .S(n_182));
   FA_X1 i_92 (.A(p_3[15]), .B(p_4[15]), .CI(p_5[15]), .CO(n_185), .S(n_184));
   FA_X1 i_93 (.A(p_6[15]), .B(p_7[15]), .CI(p_8[15]), .CO(n_187), .S(n_186));
   FA_X1 i_94 (.A(p_9[15]), .B(p_10[15]), .CI(p_11[15]), .CO(n_189), .S(n_188));
   FA_X1 i_95 (.A(p_12[15]), .B(p_13[15]), .CI(p_14[15]), .CO(n_191), .S(n_190));
   FA_X1 i_96 (.A(p_15[15]), .B(n_165), .CI(n_163), .CO(n_193), .S(n_192));
   FA_X1 i_97 (.A(n_161), .B(n_159), .CI(n_157), .CO(n_195), .S(n_194));
   FA_X1 i_98 (.A(n_167), .B(n_190), .CI(n_188), .CO(n_197), .S(n_196));
   FA_X1 i_99 (.A(n_186), .B(n_184), .CI(n_182), .CO(n_199), .S(n_198));
   FA_X1 i_100 (.A(n_169), .B(n_194), .CI(n_192), .CO(n_201), .S(n_200));
   FA_X1 i_101 (.A(n_171), .B(n_173), .CI(n_198), .CO(n_203), .S(n_202));
   FA_X1 i_102 (.A(n_196), .B(n_175), .CI(n_200), .CO(n_205), .S(n_204));
   FA_X1 i_103 (.A(n_177), .B(n_202), .CI(n_204), .CO(n_207), .S(n_206));
   HA_X1 i_104 (.A(n_179), .B(n_181), .CO(n_209), .S(n_208));
   FA_X1 i_105 (.A(p_0[16]), .B(p_1[16]), .CI(p_2[16]), .CO(n_211), .S(n_210));
   FA_X1 i_106 (.A(p_3[16]), .B(p_4[16]), .CI(p_5[16]), .CO(n_213), .S(n_212));
   FA_X1 i_107 (.A(p_6[16]), .B(p_7[16]), .CI(p_8[16]), .CO(n_215), .S(n_214));
   FA_X1 i_108 (.A(p_9[16]), .B(p_10[16]), .CI(p_11[16]), .CO(n_217), .S(n_216));
   FA_X1 i_109 (.A(p_12[16]), .B(p_13[16]), .CI(p_14[16]), .CO(n_219), .S(n_218));
   FA_X1 i_110 (.A(n_191), .B(n_189), .CI(n_187), .CO(n_221), .S(n_220));
   FA_X1 i_111 (.A(n_185), .B(n_183), .CI(n_195), .CO(n_223), .S(n_222));
   FA_X1 i_112 (.A(n_193), .B(n_218), .CI(n_216), .CO(n_225), .S(n_224));
   FA_X1 i_113 (.A(n_214), .B(n_212), .CI(n_210), .CO(n_227), .S(n_226));
   FA_X1 i_114 (.A(n_222), .B(n_220), .CI(n_199), .CO(n_229), .S(n_228));
   FA_X1 i_115 (.A(n_197), .B(n_201), .CI(n_226), .CO(n_231), .S(n_230));
   FA_X1 i_116 (.A(n_224), .B(n_228), .CI(n_203), .CO(n_233), .S(n_232));
   FA_X1 i_117 (.A(n_230), .B(n_205), .CI(n_232), .CO(n_235), .S(n_234));
   HA_X1 i_118 (.A(n_207), .B(n_209), .CO(n_237), .S(n_236));
   FA_X1 i_119 (.A(p_1[17]), .B(p_2[17]), .CI(p_3[17]), .CO(n_239), .S(n_238));
   FA_X1 i_120 (.A(p_4[17]), .B(p_5[17]), .CI(p_6[17]), .CO(n_241), .S(n_240));
   FA_X1 i_121 (.A(p_7[17]), .B(p_8[17]), .CI(p_9[17]), .CO(n_243), .S(n_242));
   FA_X1 i_122 (.A(p_10[17]), .B(p_11[17]), .CI(p_12[17]), .CO(n_245), .S(n_244));
   FA_X1 i_123 (.A(p_13[17]), .B(p_14[17]), .CI(n_219), .CO(n_247), .S(n_246));
   FA_X1 i_124 (.A(n_217), .B(n_215), .CI(n_213), .CO(n_249), .S(n_248));
   FA_X1 i_125 (.A(n_211), .B(n_221), .CI(n_246), .CO(n_251), .S(n_250));
   FA_X1 i_126 (.A(n_244), .B(n_242), .CI(n_240), .CO(n_253), .S(n_252));
   FA_X1 i_127 (.A(n_238), .B(n_223), .CI(n_248), .CO(n_255), .S(n_254));
   FA_X1 i_128 (.A(n_227), .B(n_225), .CI(n_250), .CO(n_257), .S(n_256));
   FA_X1 i_129 (.A(n_229), .B(n_252), .CI(n_254), .CO(n_259), .S(n_258));
   FA_X1 i_130 (.A(n_256), .B(n_231), .CI(n_233), .CO(n_261), .S(n_260));
   FA_X1 i_131 (.A(n_258), .B(n_260), .CI(n_235), .CO(n_263), .S(n_262));
   FA_X1 i_132 (.A(p_2[18]), .B(p_3[18]), .CI(p_4[18]), .CO(n_265), .S(n_264));
   FA_X1 i_133 (.A(p_5[18]), .B(p_6[18]), .CI(p_7[18]), .CO(n_267), .S(n_266));
   FA_X1 i_134 (.A(p_8[18]), .B(p_9[18]), .CI(p_10[18]), .CO(n_269), .S(n_268));
   FA_X1 i_135 (.A(p_11[18]), .B(p_12[18]), .CI(p_13[18]), .CO(n_271), .S(n_270));
   FA_X1 i_136 (.A(p_14[18]), .B(n_245), .CI(n_243), .CO(n_273), .S(n_272));
   FA_X1 i_137 (.A(n_241), .B(n_239), .CI(n_249), .CO(n_275), .S(n_274));
   FA_X1 i_138 (.A(n_247), .B(n_270), .CI(n_268), .CO(n_277), .S(n_276));
   FA_X1 i_139 (.A(n_266), .B(n_264), .CI(n_274), .CO(n_279), .S(n_278));
   FA_X1 i_140 (.A(n_272), .B(n_253), .CI(n_251), .CO(n_281), .S(n_280));
   FA_X1 i_141 (.A(n_255), .B(n_278), .CI(n_276), .CO(n_283), .S(n_282));
   FA_X1 i_142 (.A(n_257), .B(n_280), .CI(n_259), .CO(n_285), .S(n_284));
   FA_X1 i_143 (.A(n_282), .B(n_261), .CI(n_284), .CO(n_287), .S(n_286));
   FA_X1 i_144 (.A(p_3[19]), .B(p_4[19]), .CI(p_5[19]), .CO(n_289), .S(n_288));
   FA_X1 i_145 (.A(p_6[19]), .B(p_7[19]), .CI(p_8[19]), .CO(n_291), .S(n_290));
   FA_X1 i_146 (.A(p_9[19]), .B(p_10[19]), .CI(p_11[19]), .CO(n_293), .S(n_292));
   FA_X1 i_147 (.A(p_12[19]), .B(p_13[19]), .CI(p_14[19]), .CO(n_295), .S(n_294));
   FA_X1 i_148 (.A(n_271), .B(n_269), .CI(n_267), .CO(n_297), .S(n_296));
   FA_X1 i_149 (.A(n_265), .B(n_273), .CI(n_294), .CO(n_299), .S(n_298));
   FA_X1 i_150 (.A(n_292), .B(n_290), .CI(n_288), .CO(n_301), .S(n_300));
   FA_X1 i_151 (.A(n_275), .B(n_296), .CI(n_277), .CO(n_303), .S(n_302));
   FA_X1 i_152 (.A(n_298), .B(n_281), .CI(n_279), .CO(n_305), .S(n_304));
   FA_X1 i_153 (.A(n_300), .B(n_302), .CI(n_283), .CO(n_307), .S(n_306));
   FA_X1 i_154 (.A(n_304), .B(n_285), .CI(n_306), .CO(n_309), .S(n_308));
   FA_X1 i_155 (.A(p_4[20]), .B(p_5[20]), .CI(p_6[20]), .CO(n_311), .S(n_310));
   FA_X1 i_156 (.A(p_7[20]), .B(p_8[20]), .CI(p_9[20]), .CO(n_313), .S(n_312));
   FA_X1 i_157 (.A(p_10[20]), .B(p_11[20]), .CI(p_12[20]), .CO(n_315), .S(n_314));
   FA_X1 i_158 (.A(p_13[20]), .B(p_14[20]), .CI(n_295), .CO(n_317), .S(n_316));
   FA_X1 i_159 (.A(n_293), .B(n_291), .CI(n_289), .CO(n_319), .S(n_318));
   FA_X1 i_160 (.A(n_297), .B(n_316), .CI(n_314), .CO(n_321), .S(n_320));
   FA_X1 i_161 (.A(n_312), .B(n_310), .CI(n_318), .CO(n_323), .S(n_322));
   FA_X1 i_162 (.A(n_301), .B(n_299), .CI(n_303), .CO(n_325), .S(n_324));
   FA_X1 i_163 (.A(n_322), .B(n_320), .CI(n_305), .CO(n_327), .S(n_326));
   FA_X1 i_164 (.A(n_324), .B(n_307), .CI(n_326), .CO(n_329), .S(n_328));
   FA_X1 i_165 (.A(p_5[21]), .B(p_6[21]), .CI(p_7[21]), .CO(n_331), .S(n_330));
   FA_X1 i_166 (.A(p_8[21]), .B(p_9[21]), .CI(p_10[21]), .CO(n_333), .S(n_332));
   FA_X1 i_167 (.A(p_11[21]), .B(p_12[21]), .CI(p_13[21]), .CO(n_335), .S(n_334));
   FA_X1 i_168 (.A(p_14[21]), .B(n_315), .CI(n_313), .CO(n_337), .S(n_336));
   FA_X1 i_169 (.A(n_311), .B(n_319), .CI(n_317), .CO(n_339), .S(n_338));
   FA_X1 i_170 (.A(n_334), .B(n_332), .CI(n_330), .CO(n_341), .S(n_340));
   FA_X1 i_171 (.A(n_336), .B(n_321), .CI(n_338), .CO(n_343), .S(n_342));
   FA_X1 i_172 (.A(n_323), .B(n_340), .CI(n_325), .CO(n_345), .S(n_344));
   FA_X1 i_173 (.A(n_342), .B(n_327), .CI(n_344), .CO(n_347), .S(n_346));
   FA_X1 i_174 (.A(p_6[22]), .B(p_7[22]), .CI(p_8[22]), .CO(n_349), .S(n_348));
   FA_X1 i_175 (.A(p_9[22]), .B(p_10[22]), .CI(p_11[22]), .CO(n_351), .S(n_350));
   FA_X1 i_176 (.A(p_12[22]), .B(p_13[22]), .CI(p_14[22]), .CO(n_353), .S(n_352));
   FA_X1 i_177 (.A(n_335), .B(n_333), .CI(n_331), .CO(n_355), .S(n_354));
   FA_X1 i_178 (.A(n_337), .B(n_352), .CI(n_350), .CO(n_357), .S(n_356));
   FA_X1 i_179 (.A(n_348), .B(n_339), .CI(n_354), .CO(n_359), .S(n_358));
   FA_X1 i_180 (.A(n_341), .B(n_356), .CI(n_358), .CO(n_361), .S(n_360));
   FA_X1 i_181 (.A(n_343), .B(n_345), .CI(n_360), .CO(n_363), .S(n_362));
   FA_X1 i_182 (.A(p_7[23]), .B(p_8[23]), .CI(p_9[23]), .CO(n_365), .S(n_364));
   FA_X1 i_183 (.A(p_10[23]), .B(p_11[23]), .CI(p_12[23]), .CO(n_367), .S(n_366));
   FA_X1 i_184 (.A(p_13[23]), .B(p_14[23]), .CI(n_353), .CO(n_369), .S(n_368));
   FA_X1 i_185 (.A(n_351), .B(n_349), .CI(n_355), .CO(n_371), .S(n_370));
   FA_X1 i_186 (.A(n_368), .B(n_366), .CI(n_364), .CO(n_373), .S(n_372));
   FA_X1 i_187 (.A(n_370), .B(n_357), .CI(n_359), .CO(n_375), .S(n_374));
   FA_X1 i_188 (.A(n_372), .B(n_374), .CI(n_361), .CO(n_377), .S(n_376));
   FA_X1 i_189 (.A(p_8[24]), .B(p_9[24]), .CI(p_10[24]), .CO(n_379), .S(n_378));
   FA_X1 i_190 (.A(p_11[24]), .B(p_12[24]), .CI(p_13[24]), .CO(n_381), .S(n_380));
   FA_X1 i_191 (.A(p_14[24]), .B(n_367), .CI(n_365), .CO(n_383), .S(n_382));
   FA_X1 i_192 (.A(n_369), .B(n_380), .CI(n_378), .CO(n_385), .S(n_384));
   FA_X1 i_193 (.A(n_371), .B(n_382), .CI(n_373), .CO(n_387), .S(n_386));
   FA_X1 i_194 (.A(n_384), .B(n_375), .CI(n_386), .CO(n_389), .S(n_388));
   FA_X1 i_195 (.A(p_9[25]), .B(p_10[25]), .CI(p_11[25]), .CO(n_391), .S(n_390));
   FA_X1 i_196 (.A(p_12[25]), .B(p_13[25]), .CI(p_14[25]), .CO(n_393), .S(n_392));
   FA_X1 i_197 (.A(n_381), .B(n_379), .CI(n_383), .CO(n_395), .S(n_394));
   FA_X1 i_198 (.A(n_392), .B(n_390), .CI(n_394), .CO(n_397), .S(n_396));
   FA_X1 i_199 (.A(n_385), .B(n_387), .CI(n_396), .CO(n_399), .S(n_398));
   FA_X1 i_200 (.A(p_10[26]), .B(p_11[26]), .CI(p_12[26]), .CO(n_401), .S(n_400));
   FA_X1 i_201 (.A(p_13[26]), .B(p_14[26]), .CI(n_393), .CO(n_403), .S(n_402));
   FA_X1 i_202 (.A(n_391), .B(n_402), .CI(n_400), .CO(n_405), .S(n_404));
   FA_X1 i_203 (.A(n_395), .B(n_397), .CI(n_404), .CO(n_407), .S(n_406));
   FA_X1 i_204 (.A(p_11[27]), .B(p_12[27]), .CI(p_13[27]), .CO(n_409), .S(n_408));
   FA_X1 i_205 (.A(p_14[27]), .B(n_401), .CI(n_403), .CO(n_411), .S(n_410));
   FA_X1 i_206 (.A(n_408), .B(n_410), .CI(n_405), .CO(n_413), .S(n_412));
   FA_X1 i_207 (.A(p_12[28]), .B(p_13[28]), .CI(p_14[28]), .CO(n_415), .S(n_414));
   FA_X1 i_208 (.A(n_409), .B(n_414), .CI(n_411), .CO(n_417), .S(n_416));
   FA_X1 i_209 (.A(p_13[29]), .B(p_14[29]), .CI(n_415), .CO(n_419), .S(n_418));
   HA_X1 i_210 (.A(p_0[1]), .B(p_15[1]), .CO(n_420), .S(sum_reg[1]));
   FA_X1 i_211 (.A(p_15[2]), .B(n_0), .CI(n_420), .CO(n_421), .S(sum_reg[2]));
   FA_X1 i_212 (.A(n_4), .B(n_2), .CI(n_421), .CO(n_422), .S(sum_reg[3]));
   FA_X1 i_213 (.A(n_6), .B(n_10), .CI(n_422), .CO(n_423), .S(sum_reg[4]));
   FA_X1 i_214 (.A(n_18), .B(n_16), .CI(n_423), .CO(n_424), .S(sum_reg[5]));
   FA_X1 i_215 (.A(n_28), .B(n_26), .CI(n_424), .CO(n_425), .S(sum_reg[6]));
   FA_X1 i_216 (.A(n_38), .B(n_40), .CI(n_425), .CO(n_426), .S(sum_reg[7]));
   FA_X1 i_217 (.A(n_52), .B(n_54), .CI(n_426), .CO(n_427), .S(sum_reg[8]));
   FA_X1 i_218 (.A(n_70), .B(n_68), .CI(n_427), .CO(n_428), .S(sum_reg[9]));
   FA_X1 i_219 (.A(n_88), .B(n_86), .CI(n_428), .CO(n_429), .S(sum_reg[10]));
   FA_X1 i_220 (.A(n_106), .B(n_108), .CI(n_429), .CO(n_430), .S(sum_reg[11]));
   FA_X1 i_221 (.A(n_128), .B(n_130), .CI(n_430), .CO(n_431), .S(sum_reg[12]));
   FA_X1 i_222 (.A(n_152), .B(n_154), .CI(n_431), .CO(n_432), .S(sum_reg[13]));
   FA_X1 i_223 (.A(n_178), .B(n_180), .CI(n_432), .CO(n_433), .S(sum_reg[14]));
   FA_X1 i_224 (.A(n_206), .B(n_208), .CI(n_433), .CO(n_434), .S(sum_reg[15]));
   FA_X1 i_225 (.A(n_234), .B(n_236), .CI(n_434), .CO(n_435), .S(sum_reg[16]));
   FA_X1 i_226 (.A(n_237), .B(n_262), .CI(n_435), .CO(n_436), .S(sum_reg[17]));
   FA_X1 i_227 (.A(n_286), .B(n_263), .CI(n_436), .CO(n_437), .S(sum_reg[18]));
   FA_X1 i_228 (.A(n_287), .B(n_308), .CI(n_437), .CO(n_438), .S(sum_reg[19]));
   FA_X1 i_229 (.A(n_328), .B(n_309), .CI(n_438), .CO(n_439), .S(sum_reg[20]));
   FA_X1 i_230 (.A(n_329), .B(n_346), .CI(n_439), .CO(n_440), .S(sum_reg[21]));
   FA_X1 i_231 (.A(n_347), .B(n_362), .CI(n_440), .CO(n_441), .S(sum_reg[22]));
   FA_X1 i_232 (.A(n_376), .B(n_363), .CI(n_441), .CO(n_442), .S(sum_reg[23]));
   FA_X1 i_233 (.A(n_377), .B(n_388), .CI(n_442), .CO(n_443), .S(sum_reg[24]));
   FA_X1 i_234 (.A(n_398), .B(n_389), .CI(n_443), .CO(n_444), .S(sum_reg[25]));
   FA_X1 i_235 (.A(n_399), .B(n_406), .CI(n_444), .CO(n_445), .S(sum_reg[26]));
   FA_X1 i_236 (.A(n_412), .B(n_407), .CI(n_445), .CO(n_446), .S(sum_reg[27]));
   FA_X1 i_237 (.A(n_413), .B(n_416), .CI(n_446), .CO(n_447), .S(sum_reg[28]));
   FA_X1 i_238 (.A(n_418), .B(n_417), .CI(n_447), .CO(n_448), .S(sum_reg[29]));
   FA_X1 i_239 (.A(p_14[30]), .B(n_419), .CI(n_448), .CO(sum_reg[31]), .S(
      sum_reg[30]));
endmodule

module multiplyShiftAdd(A, B, Z);
   input [15:0]A;
   input [15:0]B;
   output [31:0]Z;

   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;

   datapath i_0_16 (.p_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_0_254, n_0_253, n_0_252, n_0_251, 
      n_0_250, n_0_249, n_0_248, n_0_247, n_0_246, n_0_245, n_0_244, n_0_243, 
      n_0_242, n_0_241, n_0_240, n_0_239, 1'b0}), .p_1({1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_0_238, 
      n_0_237, n_0_236, n_0_235, n_0_234, n_0_233, n_0_232, n_0_231, n_0_230, 
      n_0_229, n_0_228, n_0_227, n_0_226, n_0_225, n_0_224, n_0_223, 1'b0, 1'b0}), 
      .p_2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, n_0_222, n_0_221, n_0_220, n_0_219, n_0_218, n_0_217, n_0_216, 
      n_0_215, n_0_214, n_0_213, n_0_212, n_0_211, n_0_210, n_0_209, n_0_208, 
      n_0_207, 1'b0, 1'b0, 1'b0}), .p_3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_0_206, n_0_205, n_0_204, n_0_203, 
      n_0_202, n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, n_0_196, n_0_195, 
      n_0_194, n_0_193, n_0_192, n_0_191, 1'b0, 1'b0, 1'b0, 1'b0}), .p_4({1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_0_190, 
      n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, n_0_184, n_0_183, n_0_182, 
      n_0_181, n_0_180, n_0_179, n_0_178, n_0_177, n_0_176, n_0_175, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0}), .p_5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, n_0_169, n_0_168, 
      n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, n_0_161, n_0_160, 
      n_0_159, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_6({1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_0_158, n_0_157, n_0_156, n_0_155, 
      n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, 
      n_0_146, n_0_145, n_0_144, n_0_143, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0}), .p_7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_0_142, 
      n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, 
      n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_8({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
      n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
      n_0_111, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_9({
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_0_110, n_0_109, n_0_108, n_0_107, 
      n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, 
      n_0_98, n_0_97, n_0_96, n_0_95, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0}), .p_10({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_0_94, n_0_93, 
      n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, 
      n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_11({1'b0, 1'b0, 1'b0, 1'b0, n_0_78, 
      n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, 
      n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_12({1'b0, 1'b0, 1'b0, 
      n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, 
      n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_13({1'b0, 
      1'b0, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, 
      n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_14({1'b0, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
      n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0}), .p_15({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n_0_14, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, 
      n_0_1, n_0_0, uc_0}), .sum_reg({Z[31], Z[30], Z[29], Z[28], Z[27], Z[26], 
      Z[25], Z[24], Z[23], Z[22], Z[21], Z[20], Z[19], Z[18], Z[17], Z[16], 
      Z[15], Z[14], Z[13], Z[12], Z[11], Z[10], Z[9], Z[8], Z[7], Z[6], Z[5], 
      Z[4], Z[3], Z[2], Z[1], uc_1}));
   AND2_X1 i_0_0_0 (.A1(B[1]), .A2(A[0]), .ZN(n_0_239));
   AND2_X1 i_0_0_1 (.A1(B[1]), .A2(A[1]), .ZN(n_0_240));
   AND2_X1 i_0_0_2 (.A1(B[1]), .A2(A[2]), .ZN(n_0_241));
   AND2_X1 i_0_0_3 (.A1(B[1]), .A2(A[3]), .ZN(n_0_242));
   AND2_X1 i_0_0_4 (.A1(B[1]), .A2(A[4]), .ZN(n_0_243));
   AND2_X1 i_0_0_5 (.A1(B[1]), .A2(A[5]), .ZN(n_0_244));
   AND2_X1 i_0_0_6 (.A1(B[1]), .A2(A[6]), .ZN(n_0_245));
   AND2_X1 i_0_0_7 (.A1(B[1]), .A2(A[7]), .ZN(n_0_246));
   AND2_X1 i_0_0_8 (.A1(B[1]), .A2(A[8]), .ZN(n_0_247));
   AND2_X1 i_0_0_9 (.A1(B[1]), .A2(A[9]), .ZN(n_0_248));
   AND2_X1 i_0_0_10 (.A1(B[1]), .A2(A[10]), .ZN(n_0_249));
   AND2_X1 i_0_0_11 (.A1(B[1]), .A2(A[11]), .ZN(n_0_250));
   AND2_X1 i_0_0_12 (.A1(B[1]), .A2(A[12]), .ZN(n_0_251));
   AND2_X1 i_0_0_13 (.A1(B[1]), .A2(A[13]), .ZN(n_0_252));
   AND2_X1 i_0_0_14 (.A1(B[1]), .A2(A[14]), .ZN(n_0_253));
   AND2_X1 i_0_0_15 (.A1(B[1]), .A2(A[15]), .ZN(n_0_254));
   AND2_X1 i_0_0_16 (.A1(B[2]), .A2(A[0]), .ZN(n_0_223));
   AND2_X1 i_0_0_17 (.A1(B[2]), .A2(A[1]), .ZN(n_0_224));
   AND2_X1 i_0_0_18 (.A1(B[2]), .A2(A[2]), .ZN(n_0_225));
   AND2_X1 i_0_0_19 (.A1(B[2]), .A2(A[3]), .ZN(n_0_226));
   AND2_X1 i_0_0_20 (.A1(B[2]), .A2(A[4]), .ZN(n_0_227));
   AND2_X1 i_0_0_21 (.A1(B[2]), .A2(A[5]), .ZN(n_0_228));
   AND2_X1 i_0_0_22 (.A1(B[2]), .A2(A[6]), .ZN(n_0_229));
   AND2_X1 i_0_0_23 (.A1(B[2]), .A2(A[7]), .ZN(n_0_230));
   AND2_X1 i_0_0_24 (.A1(B[2]), .A2(A[8]), .ZN(n_0_231));
   AND2_X1 i_0_0_25 (.A1(B[2]), .A2(A[9]), .ZN(n_0_232));
   AND2_X1 i_0_0_26 (.A1(B[2]), .A2(A[10]), .ZN(n_0_233));
   AND2_X1 i_0_0_27 (.A1(B[2]), .A2(A[11]), .ZN(n_0_234));
   AND2_X1 i_0_0_28 (.A1(B[2]), .A2(A[12]), .ZN(n_0_235));
   AND2_X1 i_0_0_29 (.A1(B[2]), .A2(A[13]), .ZN(n_0_236));
   AND2_X1 i_0_0_30 (.A1(B[2]), .A2(A[14]), .ZN(n_0_237));
   AND2_X1 i_0_0_31 (.A1(B[2]), .A2(A[15]), .ZN(n_0_238));
   AND2_X1 i_0_0_32 (.A1(B[3]), .A2(A[0]), .ZN(n_0_207));
   AND2_X1 i_0_0_33 (.A1(B[3]), .A2(A[1]), .ZN(n_0_208));
   AND2_X1 i_0_0_34 (.A1(B[3]), .A2(A[2]), .ZN(n_0_209));
   AND2_X1 i_0_0_35 (.A1(B[3]), .A2(A[3]), .ZN(n_0_210));
   AND2_X1 i_0_0_36 (.A1(B[3]), .A2(A[4]), .ZN(n_0_211));
   AND2_X1 i_0_0_37 (.A1(B[3]), .A2(A[5]), .ZN(n_0_212));
   AND2_X1 i_0_0_38 (.A1(B[3]), .A2(A[6]), .ZN(n_0_213));
   AND2_X1 i_0_0_39 (.A1(B[3]), .A2(A[7]), .ZN(n_0_214));
   AND2_X1 i_0_0_40 (.A1(B[3]), .A2(A[8]), .ZN(n_0_215));
   AND2_X1 i_0_0_41 (.A1(B[3]), .A2(A[9]), .ZN(n_0_216));
   AND2_X1 i_0_0_42 (.A1(B[3]), .A2(A[10]), .ZN(n_0_217));
   AND2_X1 i_0_0_43 (.A1(B[3]), .A2(A[11]), .ZN(n_0_218));
   AND2_X1 i_0_0_44 (.A1(B[3]), .A2(A[12]), .ZN(n_0_219));
   AND2_X1 i_0_0_45 (.A1(B[3]), .A2(A[13]), .ZN(n_0_220));
   AND2_X1 i_0_0_46 (.A1(B[3]), .A2(A[14]), .ZN(n_0_221));
   AND2_X1 i_0_0_47 (.A1(B[3]), .A2(A[15]), .ZN(n_0_222));
   AND2_X1 i_0_0_48 (.A1(B[4]), .A2(A[0]), .ZN(n_0_191));
   AND2_X1 i_0_0_49 (.A1(B[4]), .A2(A[1]), .ZN(n_0_192));
   AND2_X1 i_0_0_50 (.A1(B[4]), .A2(A[2]), .ZN(n_0_193));
   AND2_X1 i_0_0_51 (.A1(B[4]), .A2(A[3]), .ZN(n_0_194));
   AND2_X1 i_0_0_52 (.A1(B[4]), .A2(A[4]), .ZN(n_0_195));
   AND2_X1 i_0_0_53 (.A1(B[4]), .A2(A[5]), .ZN(n_0_196));
   AND2_X1 i_0_0_54 (.A1(B[4]), .A2(A[6]), .ZN(n_0_197));
   AND2_X1 i_0_0_55 (.A1(B[4]), .A2(A[7]), .ZN(n_0_198));
   AND2_X1 i_0_0_56 (.A1(B[4]), .A2(A[8]), .ZN(n_0_199));
   AND2_X1 i_0_0_57 (.A1(B[4]), .A2(A[9]), .ZN(n_0_200));
   AND2_X1 i_0_0_58 (.A1(B[4]), .A2(A[10]), .ZN(n_0_201));
   AND2_X1 i_0_0_59 (.A1(B[4]), .A2(A[11]), .ZN(n_0_202));
   AND2_X1 i_0_0_60 (.A1(B[4]), .A2(A[12]), .ZN(n_0_203));
   AND2_X1 i_0_0_61 (.A1(B[4]), .A2(A[13]), .ZN(n_0_204));
   AND2_X1 i_0_0_62 (.A1(B[4]), .A2(A[14]), .ZN(n_0_205));
   AND2_X1 i_0_0_63 (.A1(B[4]), .A2(A[15]), .ZN(n_0_206));
   AND2_X1 i_0_0_64 (.A1(B[5]), .A2(A[0]), .ZN(n_0_175));
   AND2_X1 i_0_0_65 (.A1(B[5]), .A2(A[1]), .ZN(n_0_176));
   AND2_X1 i_0_0_66 (.A1(B[5]), .A2(A[2]), .ZN(n_0_177));
   AND2_X1 i_0_0_67 (.A1(B[5]), .A2(A[3]), .ZN(n_0_178));
   AND2_X1 i_0_0_68 (.A1(B[5]), .A2(A[4]), .ZN(n_0_179));
   AND2_X1 i_0_0_69 (.A1(B[5]), .A2(A[5]), .ZN(n_0_180));
   AND2_X1 i_0_0_70 (.A1(B[5]), .A2(A[6]), .ZN(n_0_181));
   AND2_X1 i_0_0_71 (.A1(B[5]), .A2(A[7]), .ZN(n_0_182));
   AND2_X1 i_0_0_72 (.A1(B[5]), .A2(A[8]), .ZN(n_0_183));
   AND2_X1 i_0_0_73 (.A1(B[5]), .A2(A[9]), .ZN(n_0_184));
   AND2_X1 i_0_0_74 (.A1(B[5]), .A2(A[10]), .ZN(n_0_185));
   AND2_X1 i_0_0_75 (.A1(B[5]), .A2(A[11]), .ZN(n_0_186));
   AND2_X1 i_0_0_76 (.A1(B[5]), .A2(A[12]), .ZN(n_0_187));
   AND2_X1 i_0_0_77 (.A1(B[5]), .A2(A[13]), .ZN(n_0_188));
   AND2_X1 i_0_0_78 (.A1(B[5]), .A2(A[14]), .ZN(n_0_189));
   AND2_X1 i_0_0_79 (.A1(B[5]), .A2(A[15]), .ZN(n_0_190));
   AND2_X1 i_0_0_80 (.A1(B[6]), .A2(A[0]), .ZN(n_0_159));
   AND2_X1 i_0_0_81 (.A1(B[6]), .A2(A[1]), .ZN(n_0_160));
   AND2_X1 i_0_0_82 (.A1(B[6]), .A2(A[2]), .ZN(n_0_161));
   AND2_X1 i_0_0_83 (.A1(B[6]), .A2(A[3]), .ZN(n_0_162));
   AND2_X1 i_0_0_84 (.A1(B[6]), .A2(A[4]), .ZN(n_0_163));
   AND2_X1 i_0_0_85 (.A1(B[6]), .A2(A[5]), .ZN(n_0_164));
   AND2_X1 i_0_0_86 (.A1(B[6]), .A2(A[6]), .ZN(n_0_165));
   AND2_X1 i_0_0_87 (.A1(B[6]), .A2(A[7]), .ZN(n_0_166));
   AND2_X1 i_0_0_88 (.A1(B[6]), .A2(A[8]), .ZN(n_0_167));
   AND2_X1 i_0_0_89 (.A1(B[6]), .A2(A[9]), .ZN(n_0_168));
   AND2_X1 i_0_0_90 (.A1(B[6]), .A2(A[10]), .ZN(n_0_169));
   AND2_X1 i_0_0_91 (.A1(B[6]), .A2(A[11]), .ZN(n_0_170));
   AND2_X1 i_0_0_92 (.A1(B[6]), .A2(A[12]), .ZN(n_0_171));
   AND2_X1 i_0_0_93 (.A1(B[6]), .A2(A[13]), .ZN(n_0_172));
   AND2_X1 i_0_0_94 (.A1(B[6]), .A2(A[14]), .ZN(n_0_173));
   AND2_X1 i_0_0_95 (.A1(B[6]), .A2(A[15]), .ZN(n_0_174));
   AND2_X1 i_0_0_96 (.A1(B[7]), .A2(A[0]), .ZN(n_0_143));
   AND2_X1 i_0_0_97 (.A1(B[7]), .A2(A[1]), .ZN(n_0_144));
   AND2_X1 i_0_0_98 (.A1(B[7]), .A2(A[2]), .ZN(n_0_145));
   AND2_X1 i_0_0_99 (.A1(B[7]), .A2(A[3]), .ZN(n_0_146));
   AND2_X1 i_0_0_100 (.A1(B[7]), .A2(A[4]), .ZN(n_0_147));
   AND2_X1 i_0_0_101 (.A1(B[7]), .A2(A[5]), .ZN(n_0_148));
   AND2_X1 i_0_0_102 (.A1(B[7]), .A2(A[6]), .ZN(n_0_149));
   AND2_X1 i_0_0_103 (.A1(B[7]), .A2(A[7]), .ZN(n_0_150));
   AND2_X1 i_0_0_104 (.A1(B[7]), .A2(A[8]), .ZN(n_0_151));
   AND2_X1 i_0_0_105 (.A1(B[7]), .A2(A[9]), .ZN(n_0_152));
   AND2_X1 i_0_0_106 (.A1(B[7]), .A2(A[10]), .ZN(n_0_153));
   AND2_X1 i_0_0_107 (.A1(B[7]), .A2(A[11]), .ZN(n_0_154));
   AND2_X1 i_0_0_108 (.A1(B[7]), .A2(A[12]), .ZN(n_0_155));
   AND2_X1 i_0_0_109 (.A1(B[7]), .A2(A[13]), .ZN(n_0_156));
   AND2_X1 i_0_0_110 (.A1(B[7]), .A2(A[14]), .ZN(n_0_157));
   AND2_X1 i_0_0_111 (.A1(B[7]), .A2(A[15]), .ZN(n_0_158));
   AND2_X1 i_0_0_112 (.A1(B[8]), .A2(A[0]), .ZN(n_0_127));
   AND2_X1 i_0_0_113 (.A1(B[8]), .A2(A[1]), .ZN(n_0_128));
   AND2_X1 i_0_0_114 (.A1(B[8]), .A2(A[2]), .ZN(n_0_129));
   AND2_X1 i_0_0_115 (.A1(B[8]), .A2(A[3]), .ZN(n_0_130));
   AND2_X1 i_0_0_116 (.A1(B[8]), .A2(A[4]), .ZN(n_0_131));
   AND2_X1 i_0_0_117 (.A1(B[8]), .A2(A[5]), .ZN(n_0_132));
   AND2_X1 i_0_0_118 (.A1(B[8]), .A2(A[6]), .ZN(n_0_133));
   AND2_X1 i_0_0_119 (.A1(B[8]), .A2(A[7]), .ZN(n_0_134));
   AND2_X1 i_0_0_120 (.A1(B[8]), .A2(A[8]), .ZN(n_0_135));
   AND2_X1 i_0_0_121 (.A1(B[8]), .A2(A[9]), .ZN(n_0_136));
   AND2_X1 i_0_0_122 (.A1(B[8]), .A2(A[10]), .ZN(n_0_137));
   AND2_X1 i_0_0_123 (.A1(B[8]), .A2(A[11]), .ZN(n_0_138));
   AND2_X1 i_0_0_124 (.A1(B[8]), .A2(A[12]), .ZN(n_0_139));
   AND2_X1 i_0_0_125 (.A1(B[8]), .A2(A[13]), .ZN(n_0_140));
   AND2_X1 i_0_0_126 (.A1(B[8]), .A2(A[14]), .ZN(n_0_141));
   AND2_X1 i_0_0_127 (.A1(B[8]), .A2(A[15]), .ZN(n_0_142));
   AND2_X1 i_0_0_128 (.A1(B[9]), .A2(A[0]), .ZN(n_0_111));
   AND2_X1 i_0_0_129 (.A1(B[9]), .A2(A[1]), .ZN(n_0_112));
   AND2_X1 i_0_0_130 (.A1(B[9]), .A2(A[2]), .ZN(n_0_113));
   AND2_X1 i_0_0_131 (.A1(B[9]), .A2(A[3]), .ZN(n_0_114));
   AND2_X1 i_0_0_132 (.A1(B[9]), .A2(A[4]), .ZN(n_0_115));
   AND2_X1 i_0_0_133 (.A1(B[9]), .A2(A[5]), .ZN(n_0_116));
   AND2_X1 i_0_0_134 (.A1(B[9]), .A2(A[6]), .ZN(n_0_117));
   AND2_X1 i_0_0_135 (.A1(B[9]), .A2(A[7]), .ZN(n_0_118));
   AND2_X1 i_0_0_136 (.A1(B[9]), .A2(A[8]), .ZN(n_0_119));
   AND2_X1 i_0_0_137 (.A1(B[9]), .A2(A[9]), .ZN(n_0_120));
   AND2_X1 i_0_0_138 (.A1(B[9]), .A2(A[10]), .ZN(n_0_121));
   AND2_X1 i_0_0_139 (.A1(B[9]), .A2(A[11]), .ZN(n_0_122));
   AND2_X1 i_0_0_140 (.A1(B[9]), .A2(A[12]), .ZN(n_0_123));
   AND2_X1 i_0_0_141 (.A1(B[9]), .A2(A[13]), .ZN(n_0_124));
   AND2_X1 i_0_0_142 (.A1(B[9]), .A2(A[14]), .ZN(n_0_125));
   AND2_X1 i_0_0_143 (.A1(B[9]), .A2(A[15]), .ZN(n_0_126));
   AND2_X1 i_0_0_144 (.A1(B[10]), .A2(A[0]), .ZN(n_0_95));
   AND2_X1 i_0_0_145 (.A1(B[10]), .A2(A[1]), .ZN(n_0_96));
   AND2_X1 i_0_0_146 (.A1(B[10]), .A2(A[2]), .ZN(n_0_97));
   AND2_X1 i_0_0_147 (.A1(B[10]), .A2(A[3]), .ZN(n_0_98));
   AND2_X1 i_0_0_148 (.A1(B[10]), .A2(A[4]), .ZN(n_0_99));
   AND2_X1 i_0_0_149 (.A1(B[10]), .A2(A[5]), .ZN(n_0_100));
   AND2_X1 i_0_0_150 (.A1(B[10]), .A2(A[6]), .ZN(n_0_101));
   AND2_X1 i_0_0_151 (.A1(B[10]), .A2(A[7]), .ZN(n_0_102));
   AND2_X1 i_0_0_152 (.A1(B[10]), .A2(A[8]), .ZN(n_0_103));
   AND2_X1 i_0_0_153 (.A1(B[10]), .A2(A[9]), .ZN(n_0_104));
   AND2_X1 i_0_0_154 (.A1(B[10]), .A2(A[10]), .ZN(n_0_105));
   AND2_X1 i_0_0_155 (.A1(B[10]), .A2(A[11]), .ZN(n_0_106));
   AND2_X1 i_0_0_156 (.A1(B[10]), .A2(A[12]), .ZN(n_0_107));
   AND2_X1 i_0_0_157 (.A1(B[10]), .A2(A[13]), .ZN(n_0_108));
   AND2_X1 i_0_0_158 (.A1(B[10]), .A2(A[14]), .ZN(n_0_109));
   AND2_X1 i_0_0_159 (.A1(B[10]), .A2(A[15]), .ZN(n_0_110));
   AND2_X1 i_0_0_160 (.A1(B[11]), .A2(A[0]), .ZN(n_0_79));
   AND2_X1 i_0_0_161 (.A1(B[11]), .A2(A[1]), .ZN(n_0_80));
   AND2_X1 i_0_0_162 (.A1(B[11]), .A2(A[2]), .ZN(n_0_81));
   AND2_X1 i_0_0_163 (.A1(B[11]), .A2(A[3]), .ZN(n_0_82));
   AND2_X1 i_0_0_164 (.A1(B[11]), .A2(A[4]), .ZN(n_0_83));
   AND2_X1 i_0_0_165 (.A1(B[11]), .A2(A[5]), .ZN(n_0_84));
   AND2_X1 i_0_0_166 (.A1(B[11]), .A2(A[6]), .ZN(n_0_85));
   AND2_X1 i_0_0_167 (.A1(B[11]), .A2(A[7]), .ZN(n_0_86));
   AND2_X1 i_0_0_168 (.A1(B[11]), .A2(A[8]), .ZN(n_0_87));
   AND2_X1 i_0_0_169 (.A1(B[11]), .A2(A[9]), .ZN(n_0_88));
   AND2_X1 i_0_0_170 (.A1(B[11]), .A2(A[10]), .ZN(n_0_89));
   AND2_X1 i_0_0_171 (.A1(B[11]), .A2(A[11]), .ZN(n_0_90));
   AND2_X1 i_0_0_172 (.A1(B[11]), .A2(A[12]), .ZN(n_0_91));
   AND2_X1 i_0_0_173 (.A1(B[11]), .A2(A[13]), .ZN(n_0_92));
   AND2_X1 i_0_0_174 (.A1(B[11]), .A2(A[14]), .ZN(n_0_93));
   AND2_X1 i_0_0_175 (.A1(B[11]), .A2(A[15]), .ZN(n_0_94));
   AND2_X1 i_0_0_176 (.A1(B[12]), .A2(A[0]), .ZN(n_0_63));
   AND2_X1 i_0_0_177 (.A1(B[12]), .A2(A[1]), .ZN(n_0_64));
   AND2_X1 i_0_0_178 (.A1(B[12]), .A2(A[2]), .ZN(n_0_65));
   AND2_X1 i_0_0_179 (.A1(B[12]), .A2(A[3]), .ZN(n_0_66));
   AND2_X1 i_0_0_180 (.A1(B[12]), .A2(A[4]), .ZN(n_0_67));
   AND2_X1 i_0_0_181 (.A1(B[12]), .A2(A[5]), .ZN(n_0_68));
   AND2_X1 i_0_0_182 (.A1(B[12]), .A2(A[6]), .ZN(n_0_69));
   AND2_X1 i_0_0_183 (.A1(B[12]), .A2(A[7]), .ZN(n_0_70));
   AND2_X1 i_0_0_184 (.A1(B[12]), .A2(A[8]), .ZN(n_0_71));
   AND2_X1 i_0_0_185 (.A1(B[12]), .A2(A[9]), .ZN(n_0_72));
   AND2_X1 i_0_0_186 (.A1(B[12]), .A2(A[10]), .ZN(n_0_73));
   AND2_X1 i_0_0_187 (.A1(B[12]), .A2(A[11]), .ZN(n_0_74));
   AND2_X1 i_0_0_188 (.A1(B[12]), .A2(A[12]), .ZN(n_0_75));
   AND2_X1 i_0_0_189 (.A1(B[12]), .A2(A[13]), .ZN(n_0_76));
   AND2_X1 i_0_0_190 (.A1(B[12]), .A2(A[14]), .ZN(n_0_77));
   AND2_X1 i_0_0_191 (.A1(B[12]), .A2(A[15]), .ZN(n_0_78));
   AND2_X1 i_0_0_192 (.A1(B[13]), .A2(A[0]), .ZN(n_0_47));
   AND2_X1 i_0_0_193 (.A1(B[13]), .A2(A[1]), .ZN(n_0_48));
   AND2_X1 i_0_0_194 (.A1(B[13]), .A2(A[2]), .ZN(n_0_49));
   AND2_X1 i_0_0_195 (.A1(B[13]), .A2(A[3]), .ZN(n_0_50));
   AND2_X1 i_0_0_196 (.A1(B[13]), .A2(A[4]), .ZN(n_0_51));
   AND2_X1 i_0_0_197 (.A1(B[13]), .A2(A[5]), .ZN(n_0_52));
   AND2_X1 i_0_0_198 (.A1(B[13]), .A2(A[6]), .ZN(n_0_53));
   AND2_X1 i_0_0_199 (.A1(B[13]), .A2(A[7]), .ZN(n_0_54));
   AND2_X1 i_0_0_200 (.A1(B[13]), .A2(A[8]), .ZN(n_0_55));
   AND2_X1 i_0_0_201 (.A1(B[13]), .A2(A[9]), .ZN(n_0_56));
   AND2_X1 i_0_0_202 (.A1(B[13]), .A2(A[10]), .ZN(n_0_57));
   AND2_X1 i_0_0_203 (.A1(B[13]), .A2(A[11]), .ZN(n_0_58));
   AND2_X1 i_0_0_204 (.A1(B[13]), .A2(A[12]), .ZN(n_0_59));
   AND2_X1 i_0_0_205 (.A1(B[13]), .A2(A[13]), .ZN(n_0_60));
   AND2_X1 i_0_0_206 (.A1(B[13]), .A2(A[14]), .ZN(n_0_61));
   AND2_X1 i_0_0_207 (.A1(B[13]), .A2(A[15]), .ZN(n_0_62));
   AND2_X1 i_0_0_208 (.A1(B[14]), .A2(A[0]), .ZN(n_0_31));
   AND2_X1 i_0_0_209 (.A1(B[14]), .A2(A[1]), .ZN(n_0_32));
   AND2_X1 i_0_0_210 (.A1(B[14]), .A2(A[2]), .ZN(n_0_33));
   AND2_X1 i_0_0_211 (.A1(B[14]), .A2(A[3]), .ZN(n_0_34));
   AND2_X1 i_0_0_212 (.A1(B[14]), .A2(A[4]), .ZN(n_0_35));
   AND2_X1 i_0_0_213 (.A1(B[14]), .A2(A[5]), .ZN(n_0_36));
   AND2_X1 i_0_0_214 (.A1(B[14]), .A2(A[6]), .ZN(n_0_37));
   AND2_X1 i_0_0_215 (.A1(B[14]), .A2(A[7]), .ZN(n_0_38));
   AND2_X1 i_0_0_216 (.A1(B[14]), .A2(A[8]), .ZN(n_0_39));
   AND2_X1 i_0_0_217 (.A1(B[14]), .A2(A[9]), .ZN(n_0_40));
   AND2_X1 i_0_0_218 (.A1(B[14]), .A2(A[10]), .ZN(n_0_41));
   AND2_X1 i_0_0_219 (.A1(B[14]), .A2(A[11]), .ZN(n_0_42));
   AND2_X1 i_0_0_220 (.A1(B[14]), .A2(A[12]), .ZN(n_0_43));
   AND2_X1 i_0_0_221 (.A1(B[14]), .A2(A[13]), .ZN(n_0_44));
   AND2_X1 i_0_0_222 (.A1(B[14]), .A2(A[14]), .ZN(n_0_45));
   AND2_X1 i_0_0_223 (.A1(B[14]), .A2(A[15]), .ZN(n_0_46));
   AND2_X1 i_0_0_224 (.A1(B[15]), .A2(A[0]), .ZN(n_0_15));
   AND2_X1 i_0_0_225 (.A1(B[15]), .A2(A[1]), .ZN(n_0_16));
   AND2_X1 i_0_0_226 (.A1(B[15]), .A2(A[2]), .ZN(n_0_17));
   AND2_X1 i_0_0_227 (.A1(B[15]), .A2(A[3]), .ZN(n_0_18));
   AND2_X1 i_0_0_228 (.A1(B[15]), .A2(A[4]), .ZN(n_0_19));
   AND2_X1 i_0_0_229 (.A1(B[15]), .A2(A[5]), .ZN(n_0_20));
   AND2_X1 i_0_0_230 (.A1(B[15]), .A2(A[6]), .ZN(n_0_21));
   AND2_X1 i_0_0_231 (.A1(B[15]), .A2(A[7]), .ZN(n_0_22));
   AND2_X1 i_0_0_232 (.A1(B[15]), .A2(A[8]), .ZN(n_0_23));
   AND2_X1 i_0_0_233 (.A1(B[15]), .A2(A[9]), .ZN(n_0_24));
   AND2_X1 i_0_0_234 (.A1(B[15]), .A2(A[10]), .ZN(n_0_25));
   AND2_X1 i_0_0_235 (.A1(B[15]), .A2(A[11]), .ZN(n_0_26));
   AND2_X1 i_0_0_236 (.A1(B[15]), .A2(A[12]), .ZN(n_0_27));
   AND2_X1 i_0_0_237 (.A1(B[15]), .A2(A[13]), .ZN(n_0_28));
   AND2_X1 i_0_0_238 (.A1(B[15]), .A2(A[14]), .ZN(n_0_29));
   AND2_X1 i_0_0_239 (.A1(B[15]), .A2(A[15]), .ZN(n_0_30));
   AND2_X1 i_0_0_240 (.A1(B[0]), .A2(A[0]), .ZN(Z[0]));
   AND2_X1 i_0_0_241 (.A1(B[0]), .A2(A[1]), .ZN(n_0_0));
   AND2_X1 i_0_0_242 (.A1(B[0]), .A2(A[2]), .ZN(n_0_1));
   AND2_X1 i_0_0_243 (.A1(B[0]), .A2(A[3]), .ZN(n_0_2));
   AND2_X1 i_0_0_244 (.A1(B[0]), .A2(A[4]), .ZN(n_0_3));
   AND2_X1 i_0_0_245 (.A1(B[0]), .A2(A[5]), .ZN(n_0_4));
   AND2_X1 i_0_0_246 (.A1(B[0]), .A2(A[6]), .ZN(n_0_5));
   AND2_X1 i_0_0_247 (.A1(B[0]), .A2(A[7]), .ZN(n_0_6));
   AND2_X1 i_0_0_248 (.A1(B[0]), .A2(A[8]), .ZN(n_0_7));
   AND2_X1 i_0_0_249 (.A1(B[0]), .A2(A[9]), .ZN(n_0_8));
   AND2_X1 i_0_0_250 (.A1(B[0]), .A2(A[10]), .ZN(n_0_9));
   AND2_X1 i_0_0_251 (.A1(B[0]), .A2(A[11]), .ZN(n_0_10));
   AND2_X1 i_0_0_252 (.A1(B[0]), .A2(A[12]), .ZN(n_0_11));
   AND2_X1 i_0_0_253 (.A1(B[0]), .A2(A[13]), .ZN(n_0_12));
   AND2_X1 i_0_0_254 (.A1(B[0]), .A2(A[14]), .ZN(n_0_13));
   AND2_X1 i_0_0_255 (.A1(B[0]), .A2(A[15]), .ZN(n_0_14));
endmodule
